module router_ravenoc (clk,arst,north_send,north_recv,south_send,south_recv,west_send,west_recv,east_send,east_recv,local_send,local_recv);

	input clk;
	input arst;
	input north_send;
	input west_recv;
	input east_send;
	input east_recv;
	input north_recv;
	input south_send;
	input south_recv;
	input west_send;
	input local_send;
	input local_recv;
	
	wire south_recv_resp,south_recv_req,south_send_resp,south_send_req,west_recv_resp,west_recv_req,west_send_resp,west_send_req,north_recv_resp,north_recv_req,north_send_resp,north_send_req,east_recv_resp,east_recv_req,east_send_resp,east_send_req,local_recv_resp,local_recv_req,local_send_resp,local_send_req;
	wire [194:0] int_req_v;
	wire [4:0] int_resp_v;
	wire [24:0] int_route_v;
	wire [739:0] int_map_req_v;
	wire [19:0] int_map_resp_v;
	wire [194:0] ext_req_v_i;
	wire [4:0] ext_resp_v_o;
	wire [194:0] ext_req_v_o;
	wire [4:0] ext_resp_v_i;
	wire [11:0] valid_from_im_output_module;
	wire [11:0] grant_im_output_module;
	wire [2:0] tail_flit_im_output_module;
	wire [1:0] vc_ch_act_out_output_module;
	wire req_out_output_module,xnor1resu1_output_module,xnor2resu1_output_module,and1resu1_output_module,xor1resu1_output_module,and2resu1_output_module,head_flit_output_module_32_not_output_module,and3resu1_output_module,nor23resu1_output_module,nor23resu2_output_module,and4resu1_output_module,and5resu1_output_module,or12resu12_output_module,nor23resu3_output_module,and6resu1_output_module,nand1resu_output_module,and8resu1_output_module,norfinresu1_output_module,and9resu1_output_module,and10resu1_output_module,and11resu1_output_module;
	wire [33:0] head_flit_output_module;
	wire [1:0] _sv2v_jump_output_module;
	wire [31:0] in_mod_output_module;
	wire [31:0] vc_channel_output_module;
	wire [1:0] _sv2v_jump_output_module_1;
	wire [31:0] i_output_module;
    wire [1:0] mask_ff_rr_arbiter, next_mask_rr_arbiter, mask_req_rr_arbiter, _sv2v_jump_rr_rr_arbiter, i_rr_arbiter, j_rr_arbiter, raw_grant_rr_arbiter, masked_grant_rr_arbiter, temp_mask_ff_rr_arbiter, _sv2v_jump_high_prior_arbiter1, i_high_prior_arbiter1, _sv2v_jump_high_prior_arbiter2, i_high_prior_arbiter2, mask_ff_rr_arbiter1, next_mask_rr_arbiter1, mask_req_rr_arbiter1, _sv2v_jump_rr_rr_arbiter1, i_rr_arbiter1, j_rr_arbiter1, raw_grant_rr_arbiter1, masked_grant_rr_arbiter1, temp_mask_ff_rr_arbiter11, _sv2v_jump_high_prior_arbiter11, i_high_prior_arbiter11, _sv2v_jump_high_prior_arbiter21, i_high_prior_arbiter21,mask_ff_rr_arbiter2,next_mask_rr_arbiter2,mask_req_rr_arbiter2,_sv2v_jump_rr_rr_arbiter2,i_rr_arbiter2,j_rr_arbiter2,raw_grant_rr_arbiter2,masked_grant_rr_arbiter2,temp_mask_ff_rr_arbiter22,_sv2v_jump_high_prior_arbiter12,i_high_prior_arbiter12,_sv2v_jump_high_prior_arbiter22,i_high_prior_arbiter22;

    wire xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter,xnor1res_rr_arbiter,firstif_rr_arbiter,secondif_rr_arbiter,thirdif_rr_arbiter,fourthif_rr_arbiter,not_i_rr_arbiter,arst_value_rr_arbiter,xnores_high_prior_arbiter1,i_0_not_high_prior_arbiter1,nandres_high_prior_arbiter1,xnores_high_prior_arbiter2,i_0_not_high_prior_arbiter2,nandres_high_prior_arbiter2,xnor0res_rr_arbiter1,xnor1res_rr_arbiter1,firstif_rr_arbiter1,secondif_rr_arbiter1,thirdif_rr_arbiter1,fourthif_rr_arbiter1,not_i_rr_arbiter11,arst_value_rr_arbiter1,xnores_high_prior_arbiter11,i_0_not_high_prior_arbiter11,nandres_high_prior_arbiter11,xnores_high_prior_arbiter22,i_0_not_high_prior_arbiter22,nandres_high_prior_arbiter22,xnor0res_rr_arbiter2,xnor1res_rr_arbiter2,firstif_rr_arbiter2,secondif_rr_arbiter2,thirdif_rr_arbiter2,fourthif_rr_arbiter2,not_i_rr_arbiter22,arst_value_rr_arbiter2,xnores_high_prior_arbiter12,i_0_not_high_prior_arbiter12,nandres_high_prior_arbiter12;

    wire [11:0] valid_from_im_output_module1;
    wire [11:0] grant_im_output_module1;
    wire [2:0] tail_flit_im_output_module1;
    wire [1:0] vc_ch_act_out_output_module1;
    wire req_out_output_module1,xnor1resu1_output_module1,xnor2resu1_output_module1,and1resu1_output_module1,xor1resu1_output_module1,and2resu1_output_module1,head_flit_output_module1_32_not_output_module1,and3resu1_output_module1,nor23resu1_output_module1,nor23resu2_output_module1,and4resu1_output_module1,and5resu1_output_module1,or12resu12_output_module1,nor23resu3_output_module1,and6resu1_output_module1,nand1resu_output_module1,and8resu1_output_module1,norfinresu1_output_module1,and9resu1_output_module1,and10resu1_output_module1,and11resu1_output_module1;
    wire [33:0] head_flit_output_module1;
    wire [1:0] _sv2v_jump_output_module1;
    wire [31:0] in_mod_output_module1;
    wire [31:0] vc_channel_output_module1;
    wire [1:0] _sv2v_jump_output_module1_1;
    wire [31:0] i_output_module1;
    wire [1:0] mask_ff_rr_arbiter11, next_mask_rr_arbiter11, mask_req_rr_arbiter11, _sv2v_jump_rr_rr_arbiter11, i_rr_arbiter11, j_rr_arbiter11, raw_grant_rr_arbiter11, masked_grant_rr_arbiter11, temp_mask_ff_rr_arbiter1111, _sv2v_jump_high_prior_arbiter111, i_high_prior_arbiter111, _sv2v_jump_high_prior_arbiter211, i_high_prior_arbiter211, mask_ff_rr_arbiter111, next_mask_rr_arbiter111, mask_req_rr_arbiter111, _sv2v_jump_rr_rr_arbiter111, i_rr_arbiter111, j_rr_arbiter111, raw_grant_rr_arbiter111, masked_grant_rr_arbiter111, temp_mask_ff_rr_arbiter111111, _sv2v_jump_high_prior_arbiter1111, i_high_prior_arbiter1111, _sv2v_jump_high_prior_arbiter2111, i_high_prior_arbiter2111,mask_ff_rr_arbiter112,next_mask_rr_arbiter112,mask_req_rr_arbiter112,_sv2v_jump_rr_rr_arbiter112,i_rr_arbiter112,j_rr_arbiter112,raw_grant_rr_arbiter112,masked_grant_rr_arbiter112,temp_mask_ff_rr_arbiter111122,_sv2v_jump_high_prior_arbiter1112,i_high_prior_arbiter1112,_sv2v_jump_high_prior_arbiter2112,i_high_prior_arbiter2112;

    wire xnores_high_prior_arbiter2111,i_0_not_high_prior_arbiter2111,nandres_high_prior_arbiter2111,xnor0res_rr_arbiter11,xnor1res_rr_arbiter11,firstif_rr_arbiter11,secondif_rr_arbiter11,thirdif_rr_arbiter11,fourthif_rr_arbiter11,not_i_rr_arbiter1111,arst_value_rr_arbiter11,xnores_high_prior_arbiter111,i_0_not_high_prior_arbiter111,nandres_high_prior_arbiter111,xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter111,xnor1res_rr_arbiter111,firstif_rr_arbiter111,secondif_rr_arbiter111,thirdif_rr_arbiter111,fourthif_rr_arbiter111,not_i_rr_arbiter111111,arst_value_rr_arbiter111,xnores_high_prior_arbiter1111,i_0_not_high_prior_arbiter1111,nandres_high_prior_arbiter1111,xnores_high_prior_arbiter212,i_0_not_high_prior_arbiter212,nandres_high_prior_arbiter212,xnor0res_rr_arbiter112,xnor1res_rr_arbiter112,firstif_rr_arbiter112,secondif_rr_arbiter112,thirdif_rr_arbiter112,fourthif_rr_arbiter112,not_i_rr_arbiter111122,arst_value_rr_arbiter112,xnores_high_prior_arbiter1112,i_0_not_high_prior_arbiter1112,nandres_high_prior_arbiter1112;

    wire [11:0] valid_from_im_output_module2;
    wire [11:0] grant_im_output_module2;
    wire [2:0] tail_flit_im_output_module2;
    wire [1:0] vc_ch_act_out_output_module2;
    wire req_out_output_module2,xnor1resu1_output_module2,xnor2resu1_output_module2,and1resu1_output_module2,xor1resu1_output_module2,and2resu1_output_module2,head_flit_output_module2_32_not_output_module2,and3resu1_output_module2,nor23resu1_output_module2,nor23resu2_output_module2,and4resu1_output_module2,and5resu1_output_module2,or12resu12_output_module2,nor23resu3_output_module2,and6resu1_output_module2,nand1resu_output_module2,and8resu1_output_module2,norfinresu1_output_module2,and9resu1_output_module2,and10resu1_output_module2,and11resu1_output_module2;
    wire [33:0] head_flit_output_module2;
    wire [1:0] _sv2v_jump_output_module2;
    wire [31:0] in_mod_output_module2;
    wire [31:0] vc_channel_output_module2;
    wire [1:0] _sv2v_jump_output_module2_1;
    wire [31:0] i_output_module2;
    wire [1:0] mask_ff_rr_arbiter22, next_mask_rr_arbiter22, mask_req_rr_arbiter22, _sv2v_jump_rr_rr_arbiter22, i_rr_arbiter22, j_rr_arbiter22, raw_grant_rr_arbiter22, masked_grant_rr_arbiter22, temp_mask_ff_rr_arbiter2222, _sv2v_jump_high_prior_arbiter122, i_high_prior_arbiter122, _sv2v_jump_high_prior_arbiter222, i_high_prior_arbiter222, mask_ff_rr_arbiter221, next_mask_rr_arbiter221, mask_req_rr_arbiter221, _sv2v_jump_rr_rr_arbiter221, i_rr_arbiter221, j_rr_arbiter221, raw_grant_rr_arbiter221, masked_grant_rr_arbiter221, temp_mask_ff_rr_arbiter222211, _sv2v_jump_high_prior_arbiter1221, i_high_prior_arbiter1221, _sv2v_jump_high_prior_arbiter2221, i_high_prior_arbiter2221,mask_ff_rr_arbiter222,next_mask_rr_arbiter222,mask_req_rr_arbiter222,_sv2v_jump_rr_rr_arbiter222,i_rr_arbiter222,j_rr_arbiter222,raw_grant_rr_arbiter222,masked_grant_rr_arbiter222,temp_mask_ff_rr_arbiter222222,_sv2v_jump_high_prior_arbiter1222,i_high_prior_arbiter1222,_sv2v_jump_high_prior_arbiter2222,i_high_prior_arbiter2222;

    wire xnores_high_prior_arbiter22212,i_0_not_high_prior_arbiter22212,nandres_high_prior_arbiter22212,xnor0res_rr_arbiter22,xnor1res_rr_arbiter22,firstif_rr_arbiter22,secondif_rr_arbiter22,thirdif_rr_arbiter22,fourthif_rr_arbiter22,not_i_rr_arbiter2222,arst_value_rr_arbiter22,xnores_high_prior_arbiter122,i_0_not_high_prior_arbiter122,nandres_high_prior_arbiter122,xnores_high_prior_arbiter222,i_0_not_high_prior_arbiter222,nandres_high_prior_arbiter222,xnor0res_rr_arbiter221,xnor1res_rr_arbiter221,firstif_rr_arbiter221,secondif_rr_arbiter221,thirdif_rr_arbiter221,fourthif_rr_arbiter221,not_i_rr_arbiter222211,arst_value_rr_arbiter221,xnores_high_prior_arbiter1221,i_0_not_high_prior_arbiter1221,nandres_high_prior_arbiter1221,xnores_high_prior_arbiter2222,i_0_not_high_prior_arbiter2222,nandres_high_prior_arbiter2222,xnor0res_rr_arbiter222,xnor1res_rr_arbiter222,firstif_rr_arbiter222,secondif_rr_arbiter222,thirdif_rr_arbiter222,fourthif_rr_arbiter222,not_i_rr_arbiter222222,arst_value_rr_arbiter222,xnores_high_prior_arbiter1222,i_0_not_high_prior_arbiter1222,nandres_high_prior_arbiter1222;


    wire [11:0] valid_from_im_output_module3;
    wire [11:0] grant_im_output_module3;
    wire [2:0] tail_flit_im_output_module3;
    wire [1:0] vc_ch_act_out_output_module3;
    wire req_out_output_module3,xnor1resu1_output_module3,xnor2resu1_output_module3,and1resu1_output_module3,xor1resu1_output_module3,and2resu1_output_module3,head_flit_output_module3_32_not_output_module3,and3resu1_output_module3,nor23resu1_output_module3,nor23resu2_output_module3,and4resu1_output_module3,and5resu1_output_module3,or12resu12_output_module3,nor23resu3_output_module3,and6resu1_output_module3,nand1resu_output_module3,and8resu1_output_module3,norfinresu1_output_module3,and9resu1_output_module3,and10resu1_output_module3,and11resu1_output_module3;
    wire [33:0] head_flit_output_module3;
    wire [1:0] _sv2v_jump_output_module3;
    wire [31:0] in_mod_output_module3;
    wire [31:0] vc_channel_output_module3;
    wire [1:0] _sv2v_jump_output_module3_1;
    wire [31:0] i_output_module3;
    wire [1:0] mask_ff_rr_arbiter3, next_mask_rr_arbiter3, mask_req_rr_arbiter3, _sv2v_jump_rr_rr_arbiter3, i_rr_arbiter3, j_rr_arbiter3, raw_grant_rr_arbiter3, masked_grant_rr_arbiter3, temp_mask_ff_rr_arbiter33, _sv2v_jump_high_prior_arbiter13, i_high_prior_arbiter13, _sv2v_jump_high_prior_arbiter23, i_high_prior_arbiter23, mask_ff_rr_arbiter31, next_mask_rr_arbiter31, mask_req_rr_arbiter31, _sv2v_jump_rr_rr_arbiter31, i_rr_arbiter31, j_rr_arbiter31, raw_grant_rr_arbiter31, masked_grant_rr_arbiter31, temp_mask_ff_rr_arbiter3311, _sv2v_jump_high_prior_arbiter131, i_high_prior_arbiter131, _sv2v_jump_high_prior_arbiter231, i_high_prior_arbiter231,mask_ff_rr_arbiter32,next_mask_rr_arbiter32,mask_req_rr_arbiter32,_sv2v_jump_rr_rr_arbiter32,i_rr_arbiter32,j_rr_arbiter32,raw_grant_rr_arbiter32,masked_grant_rr_arbiter32,temp_mask_ff_rr_arbiter3322,_sv2v_jump_high_prior_arbiter132,i_high_prior_arbiter132,_sv2v_jump_high_prior_arbiter232,i_high_prior_arbiter232;

    wire xnores_high_prior_arbiter2313,i_0_not_high_prior_arbiter2313,nandres_high_prior_arbiter2313,xnor0res_rr_arbiter3,xnor1res_rr_arbiter3,firstif_rr_arbiter3,secondif_rr_arbiter3,thirdif_rr_arbiter3,fourthif_rr_arbiter3,not_i_rr_arbiter33,arst_value_rr_arbiter3,xnores_high_prior_arbiter13,i_0_not_high_prior_arbiter13,nandres_high_prior_arbiter13,xnores_high_prior_arbiter23,i_0_not_high_prior_arbiter23,nandres_high_prior_arbiter23,xnor0res_rr_arbiter31,xnor1res_rr_arbiter31,firstif_rr_arbiter31,secondif_rr_arbiter31,thirdif_rr_arbiter31,fourthif_rr_arbiter31,not_i_rr_arbiter3311,arst_value_rr_arbiter31,xnores_high_prior_arbiter131,i_0_not_high_prior_arbiter131,nandres_high_prior_arbiter131,xnores_high_prior_arbiter232,i_0_not_high_prior_arbiter232,nandres_high_prior_arbiter232,xnor0res_rr_arbiter32,xnor1res_rr_arbiter32,firstif_rr_arbiter32,secondif_rr_arbiter32,thirdif_rr_arbiter32,fourthif_rr_arbiter32,not_i_rr_arbiter3322,arst_value_rr_arbiter32,xnores_high_prior_arbiter132,i_0_not_high_prior_arbiter132,nandres_high_prior_arbiter132;


    wire [11:0] valid_from_im_output_module4;
    wire [11:0] grant_im_output_module4;
    wire [2:0] tail_flit_im_output_module4;
    wire [1:0] vc_ch_act_out_output_module4;
    wire req_out_output_module4,xnor1resu1_output_module4,xnor2resu1_output_module4,and1resu1_output_module4,xor1resu1_output_module4,and2resu1_output_module4,head_flit_output_module4_32_not_output_module4,and3resu1_output_module4,nor23resu1_output_module4,nor23resu2_output_module4,and4resu1_output_module4,and5resu1_output_module4,or12resu12_output_module4,nor23resu3_output_module4,and6resu1_output_module4,nand1resu_output_module4,and8resu1_output_module4,norfinresu1_output_module4,and9resu1_output_module4,and10resu1_output_module4,and11resu1_output_module4;
    wire [33:0] head_flit_output_module4;
    wire [1:0] _sv2v_jump_output_module4;
    wire [31:0] in_mod_output_module4;
    wire [31:0] vc_channel_output_module4;
    wire [1:0] _sv2v_jump_output_module4_1;
    wire [31:0] i_output_module4;
    wire [1:0] mask_ff_rr_arbiter4, next_mask_rr_arbiter4, mask_req_rr_arbiter4, _sv2v_jump_rr_rr_arbiter4, i_rr_arbiter4, j_rr_arbiter4, raw_grant_rr_arbiter4, masked_grant_rr_arbiter4, temp_mask_ff_rr_arbiter44, _sv2v_jump_high_prior_arbiter14, i_high_prior_arbiter14, _sv2v_jump_high_prior_arbiter24, i_high_prior_arbiter24, mask_ff_rr_arbiter41, next_mask_rr_arbiter41, mask_req_rr_arbiter41, _sv2v_jump_rr_rr_arbiter41, i_rr_arbiter41, j_rr_arbiter41, raw_grant_rr_arbiter41, masked_grant_rr_arbiter41, temp_mask_ff_rr_arbiter4411, _sv2v_jump_high_prior_arbiter141, i_high_prior_arbiter141, _sv2v_jump_high_prior_arbiter241, i_high_prior_arbiter241,mask_ff_rr_arbiter42,next_mask_rr_arbiter42,mask_req_rr_arbiter42,_sv2v_jump_rr_rr_arbiter42,i_rr_arbiter42,j_rr_arbiter42,raw_grant_rr_arbiter42,masked_grant_rr_arbiter42,temp_mask_ff_rr_arbiter4422,_sv2v_jump_high_prior_arbiter142,i_high_prior_arbiter142,_sv2v_jump_high_prior_arbiter242,i_high_prior_arbiter242;

    wire xnores_high_prior_arbiter2414,i_0_not_high_prior_arbiter2414,nandres_high_prior_arbiter2414,xnor0res_rr_arbiter4,xnor1res_rr_arbiter4,firstif_rr_arbiter4,secondif_rr_arbiter4,thirdif_rr_arbiter4,fourthif_rr_arbiter4,not_i_rr_arbiter44,arst_value_rr_arbiter4,xnores_high_prior_arbiter14,i_0_not_high_prior_arbiter14,nandres_high_prior_arbiter14,xnores_high_prior_arbiter24,i_0_not_high_prior_arbiter24,nandres_high_prior_arbiter24,xnor0res_rr_arbiter41,xnor1res_rr_arbiter41,firstif_rr_arbiter41,secondif_rr_arbiter41,thirdif_rr_arbiter41,fourthif_rr_arbiter41,not_i_rr_arbiter4411,arst_value_rr_arbiter41,xnores_high_prior_arbiter141,i_0_not_high_prior_arbiter141,nandres_high_prior_arbiter141,xnores_high_prior_arbiter242,i_0_not_high_prior_arbiter242,nandres_high_prior_arbiter242,xnor0res_rr_arbiter42,xnor1res_rr_arbiter42,firstif_rr_arbiter42,secondif_rr_arbiter42,thirdif_rr_arbiter42,fourthif_rr_arbiter42,not_i_rr_arbiter4422,arst_value_rr_arbiter42,xnores_high_prior_arbiter142,i_0_not_high_prior_arbiter142,nandres_high_prior_arbiter142;

   	wire [8:0] routing_table_ff_input_router;
	wire [2:0] next_rt_input_router;
	wire [33:0] flit_input_router;
	wire new_rt_input_router,new_rt_input_routernot,norres_1_input_router,norres_2_input_router,norres_3_input_router,andfinres_input_router,and2result_input_router,norres_4_input_router,invres1_input_router,invres2_input_router,and3result_input_router,and4result_input_router,and5result_input_router,norres_5_input_router,and6result_input_router,and7result_input_router,and8result_input_router,and9result_input_router,and10result_input_router,and11result_input_router,orres1_input_router,orres2_input_router,orres3_input_router,finand1_input_router,finand2_input_router,finand3_input_router,nextrt2not_input_router,secondAndc_input_router,norres_5_input_router_2,and62result_input_router,and7result_input_router2,orres1_input_router2,finand1_input_router2,finand2_input_router2,and8result_input_router2,orres2_input_router2,and9result_input_router2,orres3_input_router2,finand3_input_router2,and11result_input_router2,nextrt2not_input_router,and10result_input_router2,arst_valuenot_input_router,finand3_input_router22;
    
    wire [8:0] routing_table_ff_input_router1;
    wire [2:0] next_rt_input_router1;
    wire [33:0] flit_input_router1;
    wire new_rt_input_router1,new_rt_input_router1not,norres_1_input_router1,norres_2_input_router1,norres_3_input_router1,andfinres_input_router1,and2result_input_router1,norres_4_input_router1,invres1_input_router1,invres2_input_router1,and3result_input_router1,and4result_input_router1,and5result_input_router1,norres_5_input_router1,and6result_input_router1,and7result_input_router1,and8result_input_router1,and9result_input_router1,and10result_input_router1,and11result_input_router1,orres1_input_router1,orres2_input_router1,orres3_input_router1,finand1_input_router1,finand2_input_router1,finand3_input_router1,nextrt2not_input_router11,secondAndc_input_router1,norres_5_input_router1_2,and62result_input_router1,and7result_input_router12,orres1_input_router12,finand1_input_router12,finand2_input_router12,and8result_input_router12,orres2_input_router12,and9result_input_router12,orres3_input_router12,finand3_input_router12,and11result_input_router12,nextrt2not_input_router11,and10result_input_router12,arst_valuenot_input_router1,finand3_input_router122;


    wire [8:0] routing_table_ff_input_router2;
    wire [2:0] next_rt_input_router2;
    wire [33:0] flit_input_router2;
    wire new_rt_input_router2,new_rt_input_router2not,norres_1_input_router2,norres_2_input_router2,norres_3_input_router2,andfinres_input_router2,and2result_input_router2,norres_4_input_router2,invres1_input_router2,invres2_input_router2,and3result_input_router2,and4result_input_router2,and5result_input_router2,norres_5_input_router2,and6result_input_router2,and7result_input_router22,and8result_input_router22,and9result_input_router22,and10result_input_router22,and11result_input_router22,orres1_input_router22,orres2_input_router22,orres3_input_router22,finand1_input_router22,finand2_input_router22,finand3_input_router222,nextrt2not_input_router22,secondAndc_input_router2,norres_5_input_router2_2,and62result_input_router2,and7result_input_router222,orres1_input_router222,finand1_input_router222,finand2_input_router222,and8result_input_router222,orres2_input_router222,and9result_input_router222,orres3_input_router222,finand3_input_router2222,and11result_input_router222,nextrt2not_input_router22,and10result_input_router222,arst_valuenot_input_router2,finand3_input_router22222;


    wire [8:0] routing_table_ff_input_router3;
    wire [2:0] next_rt_input_router3;
    wire [33:0] flit_input_router3;
    wire new_rt_input_router3,new_rt_input_router3not,norres_1_input_router3,norres_2_input_router3,norres_3_input_router3,andfinres_input_router3,and2result_input_router3,norres_4_input_router3,invres1_input_router3,invres2_input_router3,and3result_input_router3,and4result_input_router3,and5result_input_router3,norres_5_input_router3,and6result_input_router3,and7result_input_router3,and8result_input_router3,and9result_input_router3,and10result_input_router3,and11result_input_router3,orres1_input_router3,orres2_input_router3,orres3_input_router3,finand1_input_router3,finand2_input_router3,finand3_input_router3,nextrt2not_input_router33,secondAndc_input_router3,norres_5_input_router3_2,and62result_input_router3,and7result_input_router32,orres1_input_router32,finand1_input_router32,finand2_input_router32,and8result_input_router32,orres2_input_router32,and9result_input_router32,orres3_input_router32,finand3_input_router32,and11result_input_router32,nextrt2not_input_router33,and10result_input_router32,arst_valuenot_input_router3,finand3_input_router322;


    wire [8:0] routing_table_ff_input_router4;
    wire [2:0] next_rt_input_router4;
    wire [33:0] flit_input_router4;
    wire new_rt_input_router4,new_rt_input_router4not,norres_1_input_router4,norres_2_input_router4,norres_3_input_router4,andfinres_input_router4,and2result_input_router4,norres_4_input_router4,invres1_input_router4,invres2_input_router4,and3result_input_router4,and4result_input_router4,and5result_input_router4,norres_5_input_router4,and6result_input_router4,and7result_input_router4,and8result_input_router4,and9result_input_router4,and10result_input_router4,and11result_input_router4,orres1_input_router4,orres2_input_router4,orres3_input_router4,finand1_input_router4,finand2_input_router4,finand3_input_router4,nextrt2not_input_router44,secondAndc_input_router4,norres_5_input_router4_2,and62result_input_router4,and7result_input_router42,orres1_input_router42,finand1_input_router42,finand2_input_router42,and8result_input_router42,orres2_input_router42,and9result_input_router42,orres3_input_router42,finand3_input_router42,and11result_input_router42,nextrt2not_input_router44,and10result_input_router42,arst_valuenot_input_router4,finand3_input_router422;

//input router
    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router[2]) );
    BUFX1 U3(.A(flit_input_router_req_i[3]), .Y(flit_input_router[3]));
	BUFX1 U4(.A(flit_input_router_req_i[4]), .Y(flit_input_router[4]));
	BUFX1 U5(.A(flit_input_router_req_i[5]), .Y(flit_input_router[5]));
	BUFX1 U6(.A(flit_input_router_req_i[6]), .Y(flit_input_router[6]));
	BUFX1 U7(.A(flit_input_router_req_i[7]), .Y(flit_input_router[7]));
	BUFX1 U8(.A(flit_input_router_req_i[8]), .Y(flit_input_router[8]));
	BUFX1 U9(.A(flit_input_router_req_i[9]), .Y(flit_input_router[9]));
	BUFX1 U10(.A(flit_input_router_req_i[10]), .Y(flit_input_router[10]));
	BUFX1 U11(.A(flit_input_router_req_i[11]), .Y(flit_input_router[11]));
	BUFX1 U12(.A(flit_input_router_req_i[12]), .Y(flit_input_router[12]));
	BUFX1 U13(.A(flit_input_router_req_i[13]), .Y(flit_input_router[13]));
	BUFX1 U14(.A(flit_input_router_req_i[14]), .Y(flit_input_router[14]));
	BUFX1 U15(.A(flit_input_router_req_i[15]), .Y(flit_input_router[15]));
	BUFX1 U16(.A(flit_input_router_req_i[16]), .Y(flit_input_router[16]));
	BUFX1 U17(.A(flit_input_router_req_i[17]), .Y(flit_input_router[17]));
	BUFX1 U18(.A(flit_input_router_req_i[18]), .Y(flit_input_router[18]));
	BUFX1 U19(.A(flit_input_router_req_i[19]), .Y(flit_input_router[19]));
	BUFX1 U20(.A(flit_input_router_req_i[20]), .Y(flit_input_router[20]));
	BUFX1 U21(.A(flit_input_router_req_i[21]), .Y(flit_input_router[21]));
	BUFX1 U22(.A(flit_input_router_req_i[22]), .Y(flit_input_router[22]));
	BUFX1 U23(.A(flit_input_router_req_i[23]), .Y(flit_input_router[23]));
	BUFX1 U24(.A(flit_input_router_req_i[24]), .Y(flit_input_router[24]));
	BUFX1 U25(.A(flit_input_router_req_i[25]), .Y(flit_input_router[25]));
	BUFX1 U26(.A(flit_input_router_req_i[26]), .Y(flit_input_router[26]));
	BUFX1 U27(.A(flit_input_router_req_i[27]), .Y(flit_input_router[27]));
	BUFX1 U28(.A(flit_input_router_req_i[28]), .Y(flit_input_router[28]));
	BUFX1 U29(.A(flit_input_router_req_i[29]), .Y(flit_input_router[29]));
	BUFX1 U30(.A(flit_input_router_req_i[30]), .Y(flit_input_router[30]));
	BUFX1 U31(.A(flit_input_router_req_i[31]), .Y(flit_input_router[31]));
	BUFX1 U32(.A(flit_input_router_req_i[32]), .Y(flit_input_router[32]));
	BUFX1 U33(.A(flit_input_router_req_i[33]), .Y(flit_input_router[33]));
	BUFX1 U34(.A(flit_input_router_req_i[34]), .Y(flit_input_router[34]));
	BUFX1 U35(.A(flit_input_router_req_i[35]), .Y(flit_input_router[35]));
	BUFX1 U36(.A(flit_input_router_req_i[36]), .Y(flit_input_router[36]));

    NOR2X1 U37 ( .IN1(flit_input_router[33]), .IN2(flit_input_router[32]), .QN(norres_1_input_router) );
    AND2X1 U38 ( .IN1(flit_input_router_req_i[0]), .IN2(norres_1_input_router), .Q(new_rt_input_router) );

    NOR2X1 U37 ( .IN1(flit_input_router[31]), .IN2(1'b0), .QN(norres_2_input_router) );
    NOR2X1 U37 ( .IN1(flit_input_router[30]), .IN2(1'b0), .QN(norres_3_input_router) );
    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(norres_3_input_router), .Q(andfinres_input_router) );
    MUX21X1 U38 (.IN1(next_rt_input_router[0]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router[1]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router[2]), .IN2(1'b1), .S(andfinres_input_router), .Q(next_rt_input_router[2]);
    INVX1 U41 ( .A(andfinres_input_router), .Y(invres1_input_router) );


    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(invres1_input_router), .Q(and2result_input_router) );
    MUX21X1 U38 (.IN1(next_rt_input_router[0]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router[1]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router[2]), .IN2(1'b0), .S(and2result_input_router), .Q(next_rt_input_router[2]);
    INVX1 U41 ( .A(and2result_input_router), .Y(invres2_input_router) );

    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(invres1_input_router), .IN3(invres2_input_router), .Q(and3result_input_router) );
    AND2X1 U38 ( .IN1(flit_input_router[31]), .IN2(1'b1), .Q(and4result_input_router) );
    AND2X1 U38 ( .IN1(and4result_input_router), .IN2(and3result_input_router), .Q(and5result_input_router) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[2]);

   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][0]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][1]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][2]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][3]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(norres_5_input_router) );
    AND2X1 U38 ( .IN1(norres_5_input_router), .IN2(new_rt_input_router), .Q(and6result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and6result_input_router), .Q(int_route_v[4:0][4]);

    //1,2,4 and + or
    NOR2X1 U38 ( .IN1(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(and7result_input_router) );
    AND2X1 U19 ( .IN1(and7result_input_router), .IN2(next_rt_input_router[0]), .Y(orres1_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres1_input_router), .Q(finand1_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router), .Q(int_route_v[4:0][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[2]), .Q(and8result_input_router) );
    AND2X1 U19 ( .IN1(and8result_input_router), .IN2(next_rt_input_router[1]), .Y(orres2_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres2_input_router), .Q(finand2_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router), .Q(int_route_v[4:0][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and9result_input_router) );
    AND2X1 U19 ( .IN1(and9result_input_router), .IN2(next_rt_input_router[2]), .Y(orres3_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres3_input_router), .Q(finand3_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router), .Q(int_route_v[4:0][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and10result_input_router) );
    INVX1 U41 ( .A(next_rt_input_router[2]), .Y(nextrt2not_input_router) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router), .Q(and11result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    INVX1 U41 ( .A(new_rt_input_router), .Y(new_rt_input_routernot) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(flit_input_router_req_i[0]), .Q(secondAndc_input_router) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(norres_5_input_router_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router_2), .IN2(newsecondAndc_input_router_rt), .Q(and62result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and62result_input_router), .Q(int_route_v[4:0][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(and7result_input_router2) );
    AND2X1 U19 ( .IN1(and7result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .Y(orres1_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres1_input_router2), .Q(finand1_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router2), .Q(int_route_v[4:0][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Q(and8result_input_router2) );
    AND2X1 U19 ( .IN1(and8result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Y(orres2_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres2_input_router), .Q(finand2_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router2), .Q(int_route_v[4:0][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and9result_input_router2) );
    AND2X1 U19 ( .IN1(and9result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(orres3_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres3_input_router2), .Q(finand3_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router2), .Q(int_route_v[4:0][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and10result_input_router2) );
    INVX1 U41 ( .A(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(nextrt2not_input_router) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router2), .IN3(new_rt_input_routernot), .Q(and11result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(arst_valuenot_input_router), .Q(finand3_input_router22) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(next_rt_input_router[0]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(next_rt_input_router[1]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .IN2(next_rt_input_router[2]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]);    

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router1[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router1[2]) );
    BUFX1 U3(.A(flit_input_router1_req_i[3]), .Y(flit_input_router1[3]));
    BUFX1 U4(.A(flit_input_router1_req_i[4]), .Y(flit_input_router1[4]));
    BUFX1 U5(.A(flit_input_router1_req_i[5]), .Y(flit_input_router1[5]));
    BUFX1 U6(.A(flit_input_router1_req_i[6]), .Y(flit_input_router1[6]));
    BUFX1 U7(.A(flit_input_router1_req_i[7]), .Y(flit_input_router1[7]));
    BUFX1 U8(.A(flit_input_router1_req_i[8]), .Y(flit_input_router1[8]));
    BUFX1 U9(.A(flit_input_router1_req_i[9]), .Y(flit_input_router1[9]));
    BUFX1 U10(.A(flit_input_router1_req_i[10]), .Y(flit_input_router1[10]));
    BUFX1 U11(.A(flit_input_router1_req_i[11]), .Y(flit_input_router1[11]));
    BUFX1 U12(.A(flit_input_router1_req_i[12]), .Y(flit_input_router1[12]));
    BUFX1 U13(.A(flit_input_router1_req_i[13]), .Y(flit_input_router1[13]));
    BUFX1 U14(.A(flit_input_router1_req_i[14]), .Y(flit_input_router1[14]));
    BUFX1 U15(.A(flit_input_router1_req_i[15]), .Y(flit_input_router1[15]));
    BUFX1 U16(.A(flit_input_router1_req_i[16]), .Y(flit_input_router1[16]));
    BUFX1 U17(.A(flit_input_router1_req_i[17]), .Y(flit_input_router1[17]));
    BUFX1 U18(.A(flit_input_router1_req_i[18]), .Y(flit_input_router1[18]));
    BUFX1 U19(.A(flit_input_router1_req_i[19]), .Y(flit_input_router1[19]));
    BUFX1 U20(.A(flit_input_router1_req_i[20]), .Y(flit_input_router1[20]));
    BUFX1 U21(.A(flit_input_router1_req_i[21]), .Y(flit_input_router1[21]));
    BUFX1 U22(.A(flit_input_router1_req_i[22]), .Y(flit_input_router1[22]));
    BUFX1 U23(.A(flit_input_router1_req_i[23]), .Y(flit_input_router1[23]));
    BUFX1 U24(.A(flit_input_router1_req_i[24]), .Y(flit_input_router1[24]));
    BUFX1 U25(.A(flit_input_router1_req_i[25]), .Y(flit_input_router1[25]));
    BUFX1 U26(.A(flit_input_router1_req_i[26]), .Y(flit_input_router1[26]));
    BUFX1 U27(.A(flit_input_router1_req_i[27]), .Y(flit_input_router1[27]));
    BUFX1 U28(.A(flit_input_router1_req_i[28]), .Y(flit_input_router1[28]));
    BUFX1 U29(.A(flit_input_router1_req_i[29]), .Y(flit_input_router1[29]));
    BUFX1 U30(.A(flit_input_router1_req_i[30]), .Y(flit_input_router1[30]));
    BUFX1 U31(.A(flit_input_router1_req_i[31]), .Y(flit_input_router1[31]));
    BUFX1 U32(.A(flit_input_router1_req_i[32]), .Y(flit_input_router1[32]));
    BUFX1 U33(.A(flit_input_router1_req_i[33]), .Y(flit_input_router1[33]));
    BUFX1 U34(.A(flit_input_router1_req_i[34]), .Y(flit_input_router1[34]));
    BUFX1 U35(.A(flit_input_router1_req_i[35]), .Y(flit_input_router1[35]));
    BUFX1 U36(.A(flit_input_router1_req_i[36]), .Y(flit_input_router1[36]));

    NOR2X1 U37 ( .IN1(flit_input_router1[33]), .IN2(flit_input_router1[32]), .QN(norres_1_input_router1) );
    AND2X1 U38 ( .IN1(flit_input_router1_req_i[0]), .IN2(norres_1_input_router1), .Q(new_rt_input_router1) );

    NOR2X1 U37 ( .IN1(flit_input_router1[31]), .IN2(1'b0), .QN(norres_2_input_router1) );
    NOR2X1 U37 ( .IN1(flit_input_router1[30]), .IN2(1'b0), .QN(norres_3_input_router1) );
    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(norres_3_input_router1), .Q(andfinres_input_router1) );
    MUX21X1 U38 (.IN1(next_rt_input_router1[0]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[1]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[2]), .IN2(1'b1), .S(andfinres_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U41 ( .A(andfinres_input_router1), .Y(invres1_input_router1) );


    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(invres1_input_router1), .Q(and2result_input_router1) );
    MUX21X1 U38 (.IN1(next_rt_input_router1[0]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[1]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[2]), .IN2(1'b0), .S(and2result_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U41 ( .A(and2result_input_router1), .Y(invres2_input_router1) );

    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(invres1_input_router1), .IN3(invres2_input_router1), .Q(and3result_input_router1) );
    AND2X1 U38 ( .IN1(flit_input_router1[31]), .IN2(1'b1), .Q(and4result_input_router1) );
    AND2X1 U38 ( .IN1(and4result_input_router1), .IN2(and3result_input_router1), .Q(and5result_input_router1) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(norres_5_input_router1) );
    AND2X1 U38 ( .IN1(norres_5_input_router1), .IN2(new_rt_input_router1), .Q(and6result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and6result_input_router1), .Q(int_route_v[9:5][4]);

    //1,2,4 and + or
    NOR2X1 U38 ( .IN1(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(and7result_input_router1) );
    AND2X1 U19 ( .IN1(and7result_input_router1), .IN2(next_rt_input_router1[0]), .Y(orres1_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres1_input_router1), .Q(finand1_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router1), .Q(int_route_v[9:5][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[2]), .Q(and8result_input_router1) );
    AND2X1 U19 ( .IN1(and8result_input_router1), .IN2(next_rt_input_router1[1]), .Y(orres2_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres2_input_router1), .Q(finand2_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router1), .Q(int_route_v[9:5][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and9result_input_router1) );
    AND2X1 U19 ( .IN1(and9result_input_router1), .IN2(next_rt_input_router1[2]), .Y(orres3_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres3_input_router1), .Q(finand3_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router1), .Q(int_route_v[9:5][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and10result_input_router1) );
    INVX1 U41 ( .A(next_rt_input_router1[2]), .Y(nextrt2not_input_router11) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router1), .Q(and11result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    INVX1 U41 ( .A(new_rt_input_router1), .Y(new_rt_input_router1not) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(flit_input_router1_req_i[0]), .Q(secondAndc_input_router1) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(norres_5_input_router1_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router1_2), .IN2(newsecondAndc_input_router1_rt), .Q(and62result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and62result_input_router1), .Q(int_route_v[9:5][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(and7result_input_router12) );
    AND2X1 U19 ( .IN1(and7result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .Y(orres1_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres1_input_router12), .Q(finand1_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router12), .Q(int_route_v[9:5][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Q(and8result_input_router12) );
    AND2X1 U19 ( .IN1(and8result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Y(orres2_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres2_input_router1), .Q(finand2_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router12), .Q(int_route_v[9:5][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and9result_input_router12) );
    AND2X1 U19 ( .IN1(and9result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(orres3_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres3_input_router12), .Q(finand3_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router12), .Q(int_route_v[9:5][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and10result_input_router12) );
    INVX1 U41 ( .A(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(nextrt2not_input_router11) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router12), .IN3(new_rt_input_router1not), .Q(and11result_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(arst_valuenot_input_router1), .Q(finand3_input_router122) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(next_rt_input_router1[0]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(next_rt_input_router1[1]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .IN2(next_rt_input_router1[2]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]);


	BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router2[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router2[2]) );
    BUFX1 U3(.A(flit_input_router2_req_i[3]), .Y(flit_input_router2[3]));
    BUFX1 U4(.A(flit_input_router2_req_i[4]), .Y(flit_input_router2[4]));
    BUFX1 U5(.A(flit_input_router2_req_i[5]), .Y(flit_input_router2[5]));
    BUFX1 U6(.A(flit_input_router2_req_i[6]), .Y(flit_input_router2[6]));
    BUFX1 U7(.A(flit_input_router2_req_i[7]), .Y(flit_input_router2[7]));
    BUFX1 U8(.A(flit_input_router2_req_i[8]), .Y(flit_input_router2[8]));
    BUFX1 U9(.A(flit_input_router2_req_i[9]), .Y(flit_input_router2[9]));
    BUFX1 U10(.A(flit_input_router2_req_i[10]), .Y(flit_input_router2[10]));
    BUFX1 U11(.A(flit_input_router2_req_i[11]), .Y(flit_input_router2[11]));
    BUFX1 U12(.A(flit_input_router2_req_i[12]), .Y(flit_input_router2[12]));
    BUFX1 U13(.A(flit_input_router2_req_i[13]), .Y(flit_input_router2[13]));
    BUFX1 U14(.A(flit_input_router2_req_i[14]), .Y(flit_input_router2[14]));
    BUFX1 U15(.A(flit_input_router2_req_i[15]), .Y(flit_input_router2[15]));
    BUFX1 U16(.A(flit_input_router2_req_i[16]), .Y(flit_input_router2[16]));
    BUFX1 U17(.A(flit_input_router2_req_i[17]), .Y(flit_input_router2[17]));
    BUFX1 U18(.A(flit_input_router2_req_i[18]), .Y(flit_input_router2[18]));
    BUFX1 U19(.A(flit_input_router2_req_i[19]), .Y(flit_input_router2[19]));
    BUFX1 U20(.A(flit_input_router2_req_i[20]), .Y(flit_input_router2[20]));
    BUFX1 U21(.A(flit_input_router2_req_i[21]), .Y(flit_input_router2[21]));
    BUFX1 U22(.A(flit_input_router2_req_i[22]), .Y(flit_input_router2[22]));
    BUFX1 U23(.A(flit_input_router2_req_i[23]), .Y(flit_input_router2[23]));
    BUFX1 U24(.A(flit_input_router2_req_i[24]), .Y(flit_input_router2[24]));
    BUFX1 U25(.A(flit_input_router2_req_i[25]), .Y(flit_input_router2[25]));
    BUFX1 U26(.A(flit_input_router2_req_i[26]), .Y(flit_input_router2[26]));
    BUFX1 U27(.A(flit_input_router2_req_i[27]), .Y(flit_input_router2[27]));
    BUFX1 U28(.A(flit_input_router2_req_i[28]), .Y(flit_input_router2[28]));
    BUFX1 U29(.A(flit_input_router2_req_i[29]), .Y(flit_input_router2[29]));
    BUFX1 U30(.A(flit_input_router2_req_i[30]), .Y(flit_input_router2[30]));
    BUFX1 U31(.A(flit_input_router2_req_i[31]), .Y(flit_input_router2[31]));
    BUFX1 U32(.A(flit_input_router2_req_i[32]), .Y(flit_input_router2[32]));
    BUFX1 U33(.A(flit_input_router2_req_i[33]), .Y(flit_input_router2[33]));
    BUFX1 U34(.A(flit_input_router2_req_i[34]), .Y(flit_input_router2[34]));
    BUFX1 U35(.A(flit_input_router2_req_i[35]), .Y(flit_input_router2[35]));
    BUFX1 U36(.A(flit_input_router2_req_i[36]), .Y(flit_input_router2[36]));

    NOR2X1 U37 ( .IN1(flit_input_router2[33]), .IN2(flit_input_router2[32]), .QN(norres_1_input_router2) );
    AND2X1 U38 ( .IN1(flit_input_router2_req_i[0]), .IN2(norres_1_input_router2), .Q(new_rt_input_router2) );

    NOR2X1 U37 ( .IN1(flit_input_router2[31]), .IN2(1'b0), .QN(norres_2_input_router2) );
    NOR2X1 U37 ( .IN1(flit_input_router2[30]), .IN2(1'b0), .QN(norres_3_input_router2) );
    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(norres_3_input_router2), .Q(andfinres_input_router2) );
    MUX21X1 U38 (.IN1(next_rt_input_router2[0]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[1]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[2]), .IN2(1'b1), .S(andfinres_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U41 ( .A(andfinres_input_router2), .Y(invres1_input_router2) );


    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(invres1_input_router2), .Q(and2result_input_router2) );
    MUX21X1 U38 (.IN1(next_rt_input_router2[0]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[1]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[2]), .IN2(1'b0), .S(and2result_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U41 ( .A(and2result_input_router2), .Y(invres2_input_router2) );

    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(invres1_input_router2), .IN3(invres2_input_router2), .Q(and3result_input_router2) );
    AND2X1 U38 ( .IN1(flit_input_router2[31]), .IN2(1'b1), .Q(and4result_input_router2) );
    AND2X1 U38 ( .IN1(and4result_input_router2), .IN2(and3result_input_router2), .Q(and5result_input_router2) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(norres_5_input_router2) );
    AND2X1 U38 ( .IN1(norres_5_input_router2), .IN2(new_rt_input_router2), .Q(and6result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and6result_input_router2), .Q(int_route_v[14:10][4]);

    //1,2,4 and + or
    NOR2X1 U38 ( .IN1(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(and7result_input_router22) );
    AND2X1 U19 ( .IN1(and7result_input_router22), .IN2(next_rt_input_router2[0]), .Y(orres1_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres1_input_router22), .Q(finand1_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router22), .Q(int_route_v[14:10][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[2]), .Q(and8result_input_router22) );
    AND2X1 U19 ( .IN1(and8result_input_router22), .IN2(next_rt_input_router2[1]), .Y(orres2_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres2_input_router22), .Q(finand2_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router22), .Q(int_route_v[14:10][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and9result_input_router22) );
    AND2X1 U19 ( .IN1(and9result_input_router22), .IN2(next_rt_input_router2[2]), .Y(orres3_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres3_input_router22), .Q(finand3_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router222), .Q(int_route_v[14:10][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and10result_input_router22) );
    INVX1 U41 ( .A(next_rt_input_router2[2]), .Y(nextrt2not_input_router22) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router22), .Q(and11result_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    INVX1 U41 ( .A(new_rt_input_router2), .Y(new_rt_input_router2not) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(flit_input_router2_req_i[0]), .Q(secondAndc_input_router2) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(norres_5_input_router2_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router2_2), .IN2(newsecondAndc_input_router2_rt), .Q(and62result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and62result_input_router2), .Q(int_route_v[14:10][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(and7result_input_router222) );
    AND2X1 U19 ( .IN1(and7result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .Y(orres1_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres1_input_router222), .Q(finand1_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router222), .Q(int_route_v[14:10][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Q(and8result_input_router222) );
    AND2X1 U19 ( .IN1(and8result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Y(orres2_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres2_input_router22), .Q(finand2_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router222), .Q(int_route_v[14:10][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and9result_input_router222) );
    AND2X1 U19 ( .IN1(and9result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(orres3_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres3_input_router222), .Q(finand3_input_router2222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router2222), .Q(int_route_v[14:10][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and10result_input_router222) );
    INVX1 U41 ( .A(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(nextrt2not_input_router22) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router222), .IN3(new_rt_input_router2not), .Q(and11result_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(arst_valuenot_input_router2), .Q(finand3_input_router22222) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(next_rt_input_router2[0]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(next_rt_input_router2[1]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .IN2(next_rt_input_router2[2]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]); 

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router3[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router3[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router3[2]) );
    BUFX1 U3(.A(flit_input_router3_req_i[3]), .Y(flit_input_router3[3]));
    BUFX1 U4(.A(flit_input_router3_req_i[4]), .Y(flit_input_router3[4]));
    BUFX1 U5(.A(flit_input_router3_req_i[5]), .Y(flit_input_router3[5]));
    BUFX1 U6(.A(flit_input_router3_req_i[6]), .Y(flit_input_router3[6]));
    BUFX1 U7(.A(flit_input_router3_req_i[7]), .Y(flit_input_router3[7]));
    BUFX1 U8(.A(flit_input_router3_req_i[8]), .Y(flit_input_router3[8]));
    BUFX1 U9(.A(flit_input_router3_req_i[9]), .Y(flit_input_router3[9]));
    BUFX1 U10(.A(flit_input_router3_req_i[10]), .Y(flit_input_router3[10]));
    BUFX1 U11(.A(flit_input_router3_req_i[11]), .Y(flit_input_router3[11]));
    BUFX1 U12(.A(flit_input_router3_req_i[12]), .Y(flit_input_router3[12]));
    BUFX1 U13(.A(flit_input_router3_req_i[13]), .Y(flit_input_router3[13]));
    BUFX1 U14(.A(flit_input_router3_req_i[14]), .Y(flit_input_router3[14]));
    BUFX1 U15(.A(flit_input_router3_req_i[15]), .Y(flit_input_router3[15]));
    BUFX1 U16(.A(flit_input_router3_req_i[16]), .Y(flit_input_router3[16]));
    BUFX1 U17(.A(flit_input_router3_req_i[17]), .Y(flit_input_router3[17]));
    BUFX1 U18(.A(flit_input_router3_req_i[18]), .Y(flit_input_router3[18]));
    BUFX1 U19(.A(flit_input_router3_req_i[19]), .Y(flit_input_router3[19]));
    BUFX1 U20(.A(flit_input_router3_req_i[20]), .Y(flit_input_router3[20]));
    BUFX1 U21(.A(flit_input_router3_req_i[21]), .Y(flit_input_router3[21]));
    BUFX1 U22(.A(flit_input_router3_req_i[22]), .Y(flit_input_router3[22]));
    BUFX1 U23(.A(flit_input_router3_req_i[23]), .Y(flit_input_router3[23]));
    BUFX1 U24(.A(flit_input_router3_req_i[24]), .Y(flit_input_router3[24]));
    BUFX1 U25(.A(flit_input_router3_req_i[25]), .Y(flit_input_router3[25]));
    BUFX1 U26(.A(flit_input_router3_req_i[26]), .Y(flit_input_router3[26]));
    BUFX1 U27(.A(flit_input_router3_req_i[27]), .Y(flit_input_router3[27]));
    BUFX1 U28(.A(flit_input_router3_req_i[28]), .Y(flit_input_router3[28]));
    BUFX1 U29(.A(flit_input_router3_req_i[29]), .Y(flit_input_router3[29]));
    BUFX1 U30(.A(flit_input_router3_req_i[30]), .Y(flit_input_router3[30]));
    BUFX1 U31(.A(flit_input_router3_req_i[31]), .Y(flit_input_router3[31]));
    BUFX1 U32(.A(flit_input_router3_req_i[32]), .Y(flit_input_router3[32]));
    BUFX1 U33(.A(flit_input_router3_req_i[33]), .Y(flit_input_router3[33]));
    BUFX1 U34(.A(flit_input_router3_req_i[34]), .Y(flit_input_router3[34]));
    BUFX1 U35(.A(flit_input_router3_req_i[35]), .Y(flit_input_router3[35]));
    BUFX1 U36(.A(flit_input_router3_req_i[36]), .Y(flit_input_router3[36]));

    NOR2X1 U37 ( .IN1(flit_input_router3[33]), .IN2(flit_input_router3[32]), .QN(norres_1_input_router3) );
    AND2X1 U38 ( .IN1(flit_input_router3_req_i[0]), .IN2(norres_1_input_router3), .Q(new_rt_input_router3) );

    NOR2X1 U37 ( .IN1(flit_input_router3[31]), .IN2(1'b0), .QN(norres_2_input_router3) );
    NOR2X1 U37 ( .IN1(flit_input_router3[30]), .IN2(1'b0), .QN(norres_3_input_router3) );
    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(norres_3_input_router3), .Q(andfinres_input_router3) );
    MUX21X1 U38 (.IN1(next_rt_input_router3[0]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[1]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[2]), .IN2(1'b1), .S(andfinres_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U41 ( .A(andfinres_input_router3), .Y(invres1_input_router3) );


    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(invres1_input_router3), .Q(and2result_input_router3) );
    MUX21X1 U38 (.IN1(next_rt_input_router3[0]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[1]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[2]), .IN2(1'b0), .S(and2result_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U41 ( .A(and2result_input_router3), .Y(invres2_input_router3) );

    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(invres1_input_router3), .IN3(invres2_input_router3), .Q(and3result_input_router3) );
    AND2X1 U38 ( .IN1(flit_input_router3[31]), .IN2(1'b1), .Q(and4result_input_router3) );
    AND2X1 U38 ( .IN1(and4result_input_router3), .IN2(and3result_input_router3), .Q(and5result_input_router3) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(norres_5_input_router3) );
    AND2X1 U38 ( .IN1(norres_5_input_router3), .IN2(new_rt_input_router3), .Q(and6result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and6result_input_router3), .Q(int_route_v[19:15][4]);

    //1,2,4 and + or
    NOR2X1 U38 ( .IN1(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(and7result_input_router3) );
    AND2X1 U19 ( .IN1(and7result_input_router3), .IN2(next_rt_input_router3[0]), .Y(orres1_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres1_input_router3), .Q(finand1_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router3), .Q(int_route_v[19:15][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[2]), .Q(and8result_input_router3) );
    AND2X1 U19 ( .IN1(and8result_input_router3), .IN2(next_rt_input_router3[1]), .Y(orres2_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres2_input_router3), .Q(finand2_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router3), .Q(int_route_v[19:15][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and9result_input_router3) );
    AND2X1 U19 ( .IN1(and9result_input_router3), .IN2(next_rt_input_router3[2]), .Y(orres3_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres3_input_router3), .Q(finand3_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router3), .Q(int_route_v[19:15][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and10result_input_router3) );
    INVX1 U41 ( .A(next_rt_input_router3[2]), .Y(nextrt2not_input_router33) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router3), .Q(and11result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    INVX1 U41 ( .A(new_rt_input_router3), .Y(new_rt_input_router3not) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(flit_input_router3_req_i[0]), .Q(secondAndc_input_router3) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(norres_5_input_router3_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router3_2), .IN2(newsecondAndc_input_router3_rt), .Q(and62result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and62result_input_router3), .Q(int_route_v[19:15][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(and7result_input_router32) );
    AND2X1 U19 ( .IN1(and7result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .Y(orres1_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres1_input_router32), .Q(finand1_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router32), .Q(int_route_v[19:15][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Q(and8result_input_router32) );
    AND2X1 U19 ( .IN1(and8result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Y(orres2_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres2_input_router3), .Q(finand2_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router32), .Q(int_route_v[19:15][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and9result_input_router32) );
    AND2X1 U19 ( .IN1(and9result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(orres3_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres3_input_router32), .Q(finand3_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router32), .Q(int_route_v[19:15][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and10result_input_router32) );
    INVX1 U41 ( .A(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(nextrt2not_input_router33) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router32), .IN3(new_rt_input_router3not), .Q(and11result_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(arst_valuenot_input_router3), .Q(finand3_input_router322) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(next_rt_input_router3[0]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(next_rt_input_router3[1]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .IN2(next_rt_input_router3[2]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]);

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router4[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router4[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router4[2]) );
    BUFX1 U3(.A(flit_input_router4_req_i[3]), .Y(flit_input_router4[3]));
    BUFX1 U4(.A(flit_input_router4_req_i[4]), .Y(flit_input_router4[4]));
    BUFX1 U5(.A(flit_input_router4_req_i[5]), .Y(flit_input_router4[5]));
    BUFX1 U6(.A(flit_input_router4_req_i[6]), .Y(flit_input_router4[6]));
    BUFX1 U7(.A(flit_input_router4_req_i[7]), .Y(flit_input_router4[7]));
    BUFX1 U8(.A(flit_input_router4_req_i[8]), .Y(flit_input_router4[8]));
    BUFX1 U9(.A(flit_input_router4_req_i[9]), .Y(flit_input_router4[9]));
    BUFX1 U10(.A(flit_input_router4_req_i[10]), .Y(flit_input_router4[10]));
    BUFX1 U11(.A(flit_input_router4_req_i[11]), .Y(flit_input_router4[11]));
    BUFX1 U12(.A(flit_input_router4_req_i[12]), .Y(flit_input_router4[12]));
    BUFX1 U13(.A(flit_input_router4_req_i[13]), .Y(flit_input_router4[13]));
    BUFX1 U14(.A(flit_input_router4_req_i[14]), .Y(flit_input_router4[14]));
    BUFX1 U15(.A(flit_input_router4_req_i[15]), .Y(flit_input_router4[15]));
    BUFX1 U16(.A(flit_input_router4_req_i[16]), .Y(flit_input_router4[16]));
    BUFX1 U17(.A(flit_input_router4_req_i[17]), .Y(flit_input_router4[17]));
    BUFX1 U18(.A(flit_input_router4_req_i[18]), .Y(flit_input_router4[18]));
    BUFX1 U19(.A(flit_input_router4_req_i[19]), .Y(flit_input_router4[19]));
    BUFX1 U20(.A(flit_input_router4_req_i[20]), .Y(flit_input_router4[20]));
    BUFX1 U21(.A(flit_input_router4_req_i[21]), .Y(flit_input_router4[21]));
    BUFX1 U22(.A(flit_input_router4_req_i[22]), .Y(flit_input_router4[22]));
    BUFX1 U23(.A(flit_input_router4_req_i[23]), .Y(flit_input_router4[23]));
    BUFX1 U24(.A(flit_input_router4_req_i[24]), .Y(flit_input_router4[24]));
    BUFX1 U25(.A(flit_input_router4_req_i[25]), .Y(flit_input_router4[25]));
    BUFX1 U26(.A(flit_input_router4_req_i[26]), .Y(flit_input_router4[26]));
    BUFX1 U27(.A(flit_input_router4_req_i[27]), .Y(flit_input_router4[27]));
    BUFX1 U28(.A(flit_input_router4_req_i[28]), .Y(flit_input_router4[28]));
    BUFX1 U29(.A(flit_input_router4_req_i[29]), .Y(flit_input_router4[29]));
    BUFX1 U30(.A(flit_input_router4_req_i[30]), .Y(flit_input_router4[30]));
    BUFX1 U31(.A(flit_input_router4_req_i[31]), .Y(flit_input_router4[31]));
    BUFX1 U32(.A(flit_input_router4_req_i[32]), .Y(flit_input_router4[32]));
    BUFX1 U33(.A(flit_input_router4_req_i[33]), .Y(flit_input_router4[33]));
    BUFX1 U34(.A(flit_input_router4_req_i[34]), .Y(flit_input_router4[34]));
    BUFX1 U35(.A(flit_input_router4_req_i[35]), .Y(flit_input_router4[35]));
    BUFX1 U36(.A(flit_input_router4_req_i[36]), .Y(flit_input_router4[36]));

    NOR2X1 U37 ( .IN1(flit_input_router4[33]), .IN2(flit_input_router4[32]), .QN(norres_1_input_router4) );
    AND2X1 U38 ( .IN1(flit_input_router4_req_i[0]), .IN2(norres_1_input_router4), .Q(new_rt_input_router4) );

    NOR2X1 U37 ( .IN1(flit_input_router4[31]), .IN2(1'b0), .QN(norres_2_input_router4) );
    NOR2X1 U37 ( .IN1(flit_input_router4[30]), .IN2(1'b0), .QN(norres_3_input_router4) );
    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(norres_3_input_router4), .Q(andfinres_input_router4) );
    MUX21X1 U38 (.IN1(next_rt_input_router4[0]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[1]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[2]), .IN2(1'b1), .S(andfinres_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U41 ( .A(andfinres_input_router4), .Y(invres1_input_router4) );


    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(invres1_input_router4), .Q(and2result_input_router4) );
    MUX21X1 U38 (.IN1(next_rt_input_router4[0]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[1]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[2]), .IN2(1'b0), .S(and2result_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U41 ( .A(and2result_input_router4), .Y(invres2_input_router4) );

    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(invres1_input_router4), .IN3(invres2_input_router4), .Q(and3result_input_router4) );
    AND2X1 U38 ( .IN1(flit_input_router4[31]), .IN2(1'b1), .Q(and4result_input_router4) );
    AND2X1 U38 ( .IN1(and4result_input_router4), .IN2(and3result_input_router4), .Q(and5result_input_router4) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(norres_5_input_router4) );
    AND2X1 U38 ( .IN1(norres_5_input_router4), .IN2(new_rt_input_router4), .Q(and6result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and6result_input_router4), .Q(int_route_v[24:20][4]);

    //1,2,4 and + or
    NOR2X1 U38 ( .IN1(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(and7result_input_router4) );
    AND2X1 U19 ( .IN1(and7result_input_router4), .IN2(next_rt_input_router4[0]), .Y(orres1_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres1_input_router4), .Q(finand1_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router4), .Q(int_route_v[24:20][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[2]), .Q(and8result_input_router4) );
    AND2X1 U19 ( .IN1(and8result_input_router4), .IN2(next_rt_input_router4[1]), .Y(orres2_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres2_input_router4), .Q(finand2_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router4), .Q(int_route_v[24:20][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and9result_input_router4) );
    AND2X1 U19 ( .IN1(and9result_input_router4), .IN2(next_rt_input_router4[2]), .Y(orres3_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres3_input_router4), .Q(finand3_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router4), .Q(int_route_v[24:20][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and10result_input_router4) );
    INVX1 U41 ( .A(next_rt_input_router4[2]), .Y(nextrt2not_input_router44) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router4), .Q(and11result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    INVX1 U41 ( .A(new_rt_input_router4), .Y(new_rt_input_router4not) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(flit_input_router4_req_i[0]), .Q(secondAndc_input_router4) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(norres_5_input_router4_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router4_2), .IN2(newsecondAndc_input_router4_rt), .Q(and62result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and62result_input_router4), .Q(int_route_v[24:20][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(and7result_input_router42) );
    AND2X1 U19 ( .IN1(and7result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .Y(orres1_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres1_input_router42), .Q(finand1_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router42), .Q(int_route_v[24:20][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Q(and8result_input_router42) );
    AND2X1 U19 ( .IN1(and8result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Y(orres2_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres2_input_router4), .Q(finand2_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router42), .Q(int_route_v[24:20][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and9result_input_router42) );
    AND2X1 U19 ( .IN1(and9result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(orres3_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres3_input_router42), .Q(finand3_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router42), .Q(int_route_v[24:20][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and10result_input_router42) );
    INVX1 U41 ( .A(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(nextrt2not_input_router44) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router42), .IN3(new_rt_input_router4not), .Q(and11result_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(arst_valuenot_input_router4), .Q(finand3_input_router422) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(next_rt_input_router4[0]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(next_rt_input_router4[1]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .IN2(next_rt_input_router4[2]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]); 


//input part
	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[36:0]),
		.fin_resp_o(ext_resp_v_o[1:0]),
		.fout_req_o(int_req_v[36:0]),
		.fout_resp_i(int_resp_v[1:0])
	);

	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[73:37]),
		.fin_resp_o(ext_resp_v_o[2:1]),
		.fout_req_o(int_req_v[73:37]),
		.fout_resp_i(int_resp_v[2:1])
	);

	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[110:74]),
		.fin_resp_o(ext_resp_v_o[3:2]),
		.fout_req_o(int_req_v[110:74]),
		.fout_resp_i(int_resp_v[3:2])
	);

	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[147:111]),
		.fin_resp_o(ext_resp_v_o[4:3]),
		.fout_req_o(int_req_v[147:111]),
		.fout_resp_i(int_resp_v[4:3])
	);

	
	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[184:148]),
		.fin_resp_o(ext_resp_v_o[5:4]),
		.fout_req_o(int_req_v[184:148]),
		.fout_resp_i(int_resp_v[5:4])
	);


//output part	

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1[0]), .Y(i_0_not_high_prior_arbiter1) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1[0]), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(_sv2v_jump_high_prior_arbiter1[1]), .QN(nandres_high_prior_arbiter1) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2[0]), .Y(i_0_not_high_prior_arbiter2) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2[0]), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(_sv2v_jump_high_prior_arbiter2[1]), .QN(nandres_high_prior_arbiter2) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter[0]), .B(valid_from_im_output_module[3:0][0]), .Y(mask_req_rr_arbiter[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter[1]), .B(valid_from_im_output_module[3:0][1]), .Y(mask_req_rr_arbiter[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter[0]), .Y(next_mask_rr_arbiter[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter[1]), .Y(next_mask_rr_arbiter[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter[0]), .IN2(raw_grant_rr_arbiter[0]), .S(xnor0res_rr_arbiter), .Q(grant_im_output_module[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter[1]), .IN2(raw_grant_rr_arbiter[1]), .S(xnor1res_rr_arbiter), .Q(grant_im_output_module[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter[1]), .B(1'b0), .Y(firstif_rr_arbiter) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter), .B(grant_im_output_module[3:0][i_rr_arbiter[0]]), .Y(secondif_rr_arbiter) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[1]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter[0]), .Q(j_rr_arbiter[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter), .B(j_rr_arbiter[0]), .Y(thirdif_rr_arbiter) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[j_rr_arbiter[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter), .Q(next_mask_rr_arbiter[j_rr_arbiter[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b1), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(_sv2v_jump_rr_rr_arbiter[1]), .QN(fourthif_rr_arbiter) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter[0]), .IN2(next_mask_rr_arbiter[0]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter[1]), .IN2(next_mask_rr_arbiter[1]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter), .IN2(1'sb1), .S(arst_value_rr_arbiter), .Q(mask_ff_rr_arbiter[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter11) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter11[0]), .Y(i_0_not_high_prior_arbiter11) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter11), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter11[0]), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b1), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(_sv2v_jump_high_prior_arbiter11[1]), .QN(nandres_high_prior_arbiter11) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter21[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter21[0]), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(_sv2v_jump_high_prior_arbiter21[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter1[0]), .B(valid_from_im_output_module[7:4][0]), .Y(mask_req_rr_arbiter1[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter1[1]), .B(valid_from_im_output_module[7:4][1]), .Y(mask_req_rr_arbiter1[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter1[0]), .Y(next_mask_rr_arbiter1[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter1[1]), .Y(next_mask_rr_arbiter1[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter1[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter1) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter1[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter1) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter1[0]), .IN2(raw_grant_rr_arbiter1[0]), .S(xnor0res_rr_arbiter1), .Q(grant_im_output_module[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter1[1]), .IN2(raw_grant_rr_arbiter1[1]), .S(xnor1res_rr_arbiter1), .Q(grant_im_output_module[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter1[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter1[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter1[1]), .B(1'b0), .Y(firstif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter1), .B(grant_im_output_module[7:4][i_rr_arbiter1[0]]), .Y(secondif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[1]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter1[0]), .Q(j_rr_arbiter1[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter1), .B(j_rr_arbiter1[0]), .Y(thirdif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[j_rr_arbiter1[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter1), .Q(next_mask_rr_arbiter1[j_rr_arbiter1[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b1), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(_sv2v_jump_rr_rr_arbiter1[1]), .QN(fourthif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter1) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter1) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter1[0]), .IN2(next_mask_rr_arbiter1[0]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter1[1]), .IN2(next_mask_rr_arbiter1[1]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter11), .IN2(1'sb1), .S(arst_value_rr_arbiter1), .Q(mask_ff_rr_arbiter1[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter12) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter12[0]), .Y(i_0_not_high_prior_arbiter12) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter12), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter12[0]), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b1), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(_sv2v_jump_high_prior_arbiter12[1]), .QN(nandres_high_prior_arbiter12) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter22[0]), .Y(i_0_not_high_prior_arbiter22) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter22[0]), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(_sv2v_jump_high_prior_arbiter22[1]), .QN(nandres_high_prior_arbiter22) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter2[0]), .B(valid_from_im_output_module[11:8][0]), .Y(mask_req_rr_arbiter2[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter2[1]), .B(valid_from_im_output_module[11:8][1]), .Y(mask_req_rr_arbiter2[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter2[0]), .Y(next_mask_rr_arbiter2[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter2[1]), .Y(next_mask_rr_arbiter2[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter2[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter2) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter2[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter2) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter2[0]), .IN2(raw_grant_rr_arbiter2[0]), .S(xnor0res_rr_arbiter2), .Q(grant_im_output_module[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter2[1]), .IN2(raw_grant_rr_arbiter2[1]), .S(xnor1res_rr_arbiter2), .Q(grant_im_output_module[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter2[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter2[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter2[1]), .B(1'b0), .Y(firstif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter2), .B(grant_im_output_module[11:8][i_rr_arbiter2[0]]), .Y(secondif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[1]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter2[0]), .Q(j_rr_arbiter2[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter2), .B(j_rr_arbiter2[0]), .Y(thirdif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[j_rr_arbiter2[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter2), .Q(next_mask_rr_arbiter2[j_rr_arbiter2[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b1), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(_sv2v_jump_rr_rr_arbiter2[1]), .QN(fourthif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter2) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter2) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter2[0]), .IN2(next_mask_rr_arbiter2[0]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter2[1]), .IN2(next_mask_rr_arbiter2[1]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter22), .IN2(1'sb1), .S(arst_value_rr_arbiter2), .Q(mask_ff_rr_arbiter2[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37]), .IN2(vc_channel_output_module[1]), .QN(xnor1resu1_output_module) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37-1]), .IN2(vc_channel_output_module[0]), .QN(xnor2resu1_output_module) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module), .IN2(xnor2resu1_output_module), .Q(and1resu1_output_module) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]), .IN2(1'b1), .S(and1resu1_output_module), .Q(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .Q(xor1resu1_output_module) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module_1[0]), .IN2(_sv2v_jump_output_module[0]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module_1[1]), .IN2(_sv2v_jump_output_module[1]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[vc_channel_output_module[1:0]*4+in_mod_output_module[1:0]]), .Q(and2resu1_output_module) );

    MUX21X1 U3(.IN1(head_flit_output_module[3]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+3]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[3]));
	MUX21X1 U4(.IN1(head_flit_output_module[4]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+4]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[4]));
	MUX21X1 U5(.IN1(head_flit_output_module[5]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+5]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[5]));
	MUX21X1 U6(.IN1(head_flit_output_module[6]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+6]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[6]));
	MUX21X1 U7(.IN1(head_flit_output_module[7]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+7]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[7]));
	MUX21X1 U8(.IN1(head_flit_output_module[8]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+8]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[8]));
	MUX21X1 U9(.IN1(head_flit_output_module[9]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+9]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[9]));
	MUX21X1 U10(.IN1(head_flit_output_module[10]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+10]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[10]));
	MUX21X1 U11(.IN1(head_flit_output_module[11]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+11]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[11]));
	MUX21X1 U12(.IN1(head_flit_output_module[12]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+12]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[12]));
	MUX21X1 U13(.IN1(head_flit_output_module[13]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+13]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[13]));
	MUX21X1 U14(.IN1(head_flit_output_module[14]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+14]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[14]));
	MUX21X1 U15(.IN1(head_flit_output_module[15]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+15]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[15]));
	MUX21X1 U16(.IN1(head_flit_output_module[16]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+16]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[16]));
	MUX21X1 U17(.IN1(head_flit_output_module[17]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+17]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[17]));
	MUX21X1 U18(.IN1(head_flit_output_module[18]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+18]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[18]));
	MUX21X1 U19(.IN1(head_flit_output_module[19]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+19]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[19]));
	MUX21X1 U20(.IN1(head_flit_output_module[20]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+20]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[20]));
	MUX21X1 U21(.IN1(head_flit_output_module[21]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+21]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[21]));
	MUX21X1 U22(.IN1(head_flit_output_module[22]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+22]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[22]));
	MUX21X1 U23(.IN1(head_flit_output_module[23]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+23]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[23]));
	MUX21X1 U24(.IN1(head_flit_output_module[24]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+24]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[24]));
	MUX21X1 U25(.IN1(head_flit_output_module[25]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+25]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[25]));
	MUX21X1 U26(.IN1(head_flit_output_module[26]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+26]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[26]));
	MUX21X1 U27(.IN1(head_flit_output_module[27]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+27]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[27]));
	MUX21X1 U28(.IN1(head_flit_output_module[28]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+28]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[28]));
	MUX21X1 U29(.IN1(head_flit_output_module[29]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+29]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[29]));
	MUX21X1 U30(.IN1(head_flit_output_module[30]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+30]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[30]));
	MUX21X1 U31(.IN1(head_flit_output_module[31]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+31]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[31]));
	MUX21X1 U32(.IN1(head_flit_output_module[32]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+32]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[32]));
	MUX21X1 U33(.IN1(head_flit_output_module[33]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+33]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[33]));
	MUX21X1 U34(.IN1(head_flit_output_module[34]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+34]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[34]));
	MUX21X1 U35(.IN1(head_flit_output_module[35]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+35]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[35]));
	MUX21X1 U36(.IN1(head_flit_output_module[36]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+36]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[36]));

    INVX1 U041 ( .A(head_flit_output_module[32]), .Y(head_flit_output_module_32_not_output_module) );
    AND2X1 U1218 ( .IN1(head_flit_output_module_32_not_output_module), .IN2(head_flit_output_module[33]), .Q(and3resu1_output_module) );
    NOR4X1 U175821 (.IN1(head_flit_output_module[29]), .IN2(head_flit_output_module[28]), .IN3(head_flit_output_module[27]), .IN4(head_flit_output_module[26]), .Q(nor23resu1_output_module) );
    NOR4X1 U175831 (.IN1(head_flit_output_module[25]), .IN2(head_flit_output_module[24]), .IN3(head_flit_output_module[23]), .IN4(head_flit_output_module[22]), .Q(nor23resu2_output_module) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module), .IN2(nor23resu2_output_module), .Q(and4resu1_output_module) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module[33]), .IN2(head_flit_output_module[32]), .Q(nor23resu3_output_module) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module), .IN2(and4resu1_output_module), .Q(and5resu1_output_module) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module), .IN2(nor23resu3_output_module), .Q(or12resu12_output_module) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[1:0][0]), .IN2(or12resu12_output_module), .Q(and6resu1_output_module) );    
	MUX21X1 U361(.IN1(tail_flit_im_output_module[vc_channel_output_module[1:0]]), .IN2(and6resu1_output_module), .S(and2resu1_output_module) ,.Q(tail_flit_im_output_module[vc_channel_output_module[1:0]]);
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module[0]),.B(_sv2v_jump_output_module[1]),.Y(nand1resu_output_module));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module), .IN2(nand1resu_output_module), .Q(and7resu1) );    
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(_sv2v_jump_output_module_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );



	BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module[0]));
	BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[i_output_module[1:0] * 4+:4]), .Q(and8resu1_output_module) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module[0]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[0]);
	MUX21X1 U3631(.IN1(vc_ch_act_out_output_module[1]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[1]);
	MUX21X1 U3631(.IN1(req_out_output_module), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(req_out_output_module);
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module[1]), .Q(norfinresu1_output_module) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module), .IN2(req_out_output_module), .Q(and9resu1_output_module) );    
	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module), .IN2(grant_im_output_module[(vc_ch_act_out_output_module * 4) + i_output_module[1:0]]), .Q(and10resu1_output_module) );    

	MUX21X1 U3(.IN1(ext_req_v_o[36:0][3]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+3]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][3]));
	MUX21X1 U4(.IN1(ext_req_v_o[36:0][4]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+4]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][4]));
	MUX21X1 U5(.IN1(ext_req_v_o[36:0][5]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+5]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][5]));
	MUX21X1 U6(.IN1(ext_req_v_o[36:0][6]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+6]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][6]));
	MUX21X1 U7(.IN1(ext_req_v_o[36:0][7]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+7]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][7]));
	MUX21X1 U8(.IN1(ext_req_v_o[36:0][8]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+8]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][8]));
	MUX21X1 U9(.IN1(ext_req_v_o[36:0][9]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+9]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][9]));
	MUX21X1 U10(.IN1(ext_req_v_o[36:0][10]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+10]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][10]));
	MUX21X1 U11(.IN1(ext_req_v_o[36:0][11]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+11]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][11]));
	MUX21X1 U12(.IN1(ext_req_v_o[36:0][12]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+12]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][12]));
	MUX21X1 U13(.IN1(ext_req_v_o[36:0][13]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+13]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][13]));
	MUX21X1 U14(.IN1(ext_req_v_o[36:0][14]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+14]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][14]));
	MUX21X1 U15(.IN1(ext_req_v_o[36:0][15]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+15]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][15]));
	MUX21X1 U16(.IN1(ext_req_v_o[36:0][16]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+16]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][16]));
	MUX21X1 U17(.IN1(ext_req_v_o[36:0][17]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+17]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][17]));
	MUX21X1 U18(.IN1(ext_req_v_o[36:0][18]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+18]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][18]));
	MUX21X1 U19(.IN1(ext_req_v_o[36:0][19]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+19]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][19]));
	MUX21X1 U20(.IN1(ext_req_v_o[36:0][20]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+20]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][20]));
	MUX21X1 U21(.IN1(ext_req_v_o[36:0][21]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+21]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][21]));
	MUX21X1 U22(.IN1(ext_req_v_o[36:0][22]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+22]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][22]));
	MUX21X1 U23(.IN1(ext_req_v_o[36:0][23]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+23]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][23]));
	MUX21X1 U24(.IN1(ext_req_v_o[36:0][24]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+24]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][24]));
	MUX21X1 U25(.IN1(ext_req_v_o[36:0][25]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+25]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][25]));
	MUX21X1 U26(.IN1(ext_req_v_o[36:0][26]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+26]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][26]));
	MUX21X1 U27(.IN1(ext_req_v_o[36:0][27]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+27]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][27]));
	MUX21X1 U28(.IN1(ext_req_v_o[36:0][28]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+28]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][28]));
	MUX21X1 U29(.IN1(ext_req_v_o[36:0][29]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+29]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][29]));
	MUX21X1 U30(.IN1(ext_req_v_o[36:0][30]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+30]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][30]));
	MUX21X1 U31(.IN1(ext_req_v_o[36:0][31]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+31]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][31]));
	MUX21X1 U32(.IN1(ext_req_v_o[36:0][32]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+32]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][32]));
	MUX21X1 U33(.IN1(ext_req_v_o[36:0][33]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+33]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][33]));
	MUX21X1 U34(.IN1(ext_req_v_o[36:0][34]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+34]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][34]));
	MUX21X1 U35(.IN1(ext_req_v_o[36:0][35]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+35]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][35]));
	MUX21X1 U36(.IN1(ext_req_v_o[36:0][36]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+36]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][36]));

	MUX21X1 U36221(.IN1(ext_req_v_o[36:0][0]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][0]);
	MUX21X1 U36221(.IN1(ext_req_v_o[36:0][1]), .IN2(vc_ch_act_out_output_module[0]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][1]);
	MUX21X1 U36331(.IN1(ext_req_v_o[36:0][2]), .IN2(vc_ch_act_out_output_module[1]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][2]);    
	MUX21X1 U36221(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U36331(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module), .IN2(nand1resu_output_module), .Q(and11resu1_output_module) );    
	MUX21X1 U36221(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U36331(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);  





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter111[0]), .Y(i_0_not_high_prior_arbiter111) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter111), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter111[0]), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(_sv2v_jump_high_prior_arbiter111[1]), .QN(nandres_high_prior_arbiter111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter211[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter211[0]), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(_sv2v_jump_high_prior_arbiter211[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter11[0]), .B(valid_from_im_output_module1[3:0][0]), .Y(mask_req_rr_arbiter11[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter11[1]), .B(valid_from_im_output_module1[3:0][1]), .Y(mask_req_rr_arbiter11[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter11[0]), .Y(next_mask_rr_arbiter11[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter11[1]), .Y(next_mask_rr_arbiter11[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter11[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter11) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter11[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter11) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter11[0]), .IN2(raw_grant_rr_arbiter11[0]), .S(xnor0res_rr_arbiter11), .Q(grant_im_output_module1[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter11[1]), .IN2(raw_grant_rr_arbiter11[1]), .S(xnor1res_rr_arbiter11), .Q(grant_im_output_module1[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter11[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter11[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter11[1]), .B(1'b0), .Y(firstif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter11), .B(grant_im_output_module1[3:0][i_rr_arbiter11[0]]), .Y(secondif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[1]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter11[0]), .Q(j_rr_arbiter11[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter11), .B(j_rr_arbiter11[0]), .Y(thirdif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[j_rr_arbiter11[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter11), .Q(next_mask_rr_arbiter11[j_rr_arbiter11[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b1), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(_sv2v_jump_rr_rr_arbiter11[1]), .QN(fourthif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter11) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter11) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter11[0]), .IN2(next_mask_rr_arbiter11[0]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter11[1]), .IN2(next_mask_rr_arbiter11[1]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter1111), .IN2(1'sb1), .S(arst_value_rr_arbiter11), .Q(mask_ff_rr_arbiter11[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1111[0]), .Y(i_0_not_high_prior_arbiter1111) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1111), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1111[0]), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(_sv2v_jump_high_prior_arbiter1111[1]), .QN(nandres_high_prior_arbiter1111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2111[0]), .Y(i_0_not_high_prior_arbiter2111) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2111), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2111[0]), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(_sv2v_jump_high_prior_arbiter2111[1]), .QN(nandres_high_prior_arbiter2111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter111[0]), .B(valid_from_im_output_module1[7:4][0]), .Y(mask_req_rr_arbiter111[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter111[1]), .B(valid_from_im_output_module1[7:4][1]), .Y(mask_req_rr_arbiter111[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter111[0]), .Y(next_mask_rr_arbiter111[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter111[1]), .Y(next_mask_rr_arbiter111[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter111[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter111) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter111[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter111) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter111[0]), .IN2(raw_grant_rr_arbiter111[0]), .S(xnor0res_rr_arbiter111), .Q(grant_im_output_module1[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter111[1]), .IN2(raw_grant_rr_arbiter111[1]), .S(xnor1res_rr_arbiter111), .Q(grant_im_output_module1[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter111[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter111[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter111[1]), .B(1'b0), .Y(firstif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter111), .B(grant_im_output_module1[7:4][i_rr_arbiter111[0]]), .Y(secondif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[1]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter111[0]), .Q(j_rr_arbiter111[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter111), .B(j_rr_arbiter111[0]), .Y(thirdif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[j_rr_arbiter111[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter111), .Q(next_mask_rr_arbiter111[j_rr_arbiter111[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b1), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(_sv2v_jump_rr_rr_arbiter111[1]), .QN(fourthif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter111) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter111) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter111[0]), .IN2(next_mask_rr_arbiter111[0]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter111[1]), .IN2(next_mask_rr_arbiter111[1]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter111111), .IN2(1'sb1), .S(arst_value_rr_arbiter111), .Q(mask_ff_rr_arbiter111[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1112) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1112[0]), .Y(i_0_not_high_prior_arbiter1112) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1112), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1112[0]), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b1), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(_sv2v_jump_high_prior_arbiter1112[1]), .QN(nandres_high_prior_arbiter1112) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter212) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2112[0]), .Y(i_0_not_high_prior_arbiter212) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter212), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2112[0]), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(_sv2v_jump_high_prior_arbiter2112[1]), .QN(nandres_high_prior_arbiter212) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter112[0]), .B(valid_from_im_output_module1[11:8][0]), .Y(mask_req_rr_arbiter112[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter112[1]), .B(valid_from_im_output_module1[11:8][1]), .Y(mask_req_rr_arbiter112[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter112[0]), .Y(next_mask_rr_arbiter112[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter112[1]), .Y(next_mask_rr_arbiter112[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter112[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter112) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter112[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter112) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter112[0]), .IN2(raw_grant_rr_arbiter112[0]), .S(xnor0res_rr_arbiter112), .Q(grant_im_output_module1[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter112[1]), .IN2(raw_grant_rr_arbiter112[1]), .S(xnor1res_rr_arbiter112), .Q(grant_im_output_module1[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter112[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter112[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter112[1]), .B(1'b0), .Y(firstif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter112), .B(grant_im_output_module1[11:8][i_rr_arbiter112[0]]), .Y(secondif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[1]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter112[0]), .Q(j_rr_arbiter112[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter112), .B(j_rr_arbiter112[0]), .Y(thirdif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[j_rr_arbiter112[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter112), .Q(next_mask_rr_arbiter112[j_rr_arbiter112[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b1), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(_sv2v_jump_rr_rr_arbiter112[1]), .QN(fourthif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter112) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter112) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter112[0]), .IN2(next_mask_rr_arbiter112[0]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter112[1]), .IN2(next_mask_rr_arbiter112[1]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter111122), .IN2(1'sb1), .S(arst_value_rr_arbiter112), .Q(mask_ff_rr_arbiter112[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37]), .IN2(vc_channel_output_module1[1]), .QN(xnor1resu1_output_module1) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37-1]), .IN2(vc_channel_output_module1[0]), .QN(xnor2resu1_output_module1) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module1), .IN2(xnor2resu1_output_module1), .Q(and1resu1_output_module1) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]), .IN2(1'b1), .S(and1resu1_output_module1), .Q(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .Q(xor1resu1_output_module1) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module1_1[0]), .IN2(_sv2v_jump_output_module1[0]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module1_1[1]), .IN2(_sv2v_jump_output_module1[1]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[vc_channel_output_module1[1:0]*4+in_mod_output_module1[1:0]]), .Q(and2resu1_output_module1) );

    MUX21X1 U3(.IN1(head_flit_output_module1[3]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+3]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[3]));
    MUX21X1 U4(.IN1(head_flit_output_module1[4]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+4]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[4]));
    MUX21X1 U5(.IN1(head_flit_output_module1[5]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+5]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[5]));
    MUX21X1 U6(.IN1(head_flit_output_module1[6]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+6]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[6]));
    MUX21X1 U7(.IN1(head_flit_output_module1[7]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+7]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[7]));
    MUX21X1 U8(.IN1(head_flit_output_module1[8]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+8]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[8]));
    MUX21X1 U9(.IN1(head_flit_output_module1[9]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+9]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[9]));
    MUX21X1 U10(.IN1(head_flit_output_module1[10]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+10]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[10]));
    MUX21X1 U11(.IN1(head_flit_output_module1[11]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+11]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[11]));
    MUX21X1 U12(.IN1(head_flit_output_module1[12]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+12]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[12]));
    MUX21X1 U13(.IN1(head_flit_output_module1[13]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+13]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[13]));
    MUX21X1 U14(.IN1(head_flit_output_module1[14]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+14]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[14]));
    MUX21X1 U15(.IN1(head_flit_output_module1[15]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+15]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[15]));
    MUX21X1 U16(.IN1(head_flit_output_module1[16]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+16]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[16]));
    MUX21X1 U17(.IN1(head_flit_output_module1[17]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+17]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[17]));
    MUX21X1 U18(.IN1(head_flit_output_module1[18]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+18]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[18]));
    MUX21X1 U19(.IN1(head_flit_output_module1[19]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+19]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[19]));
    MUX21X1 U20(.IN1(head_flit_output_module1[20]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+20]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[20]));
    MUX21X1 U21(.IN1(head_flit_output_module1[21]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+21]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[21]));
    MUX21X1 U22(.IN1(head_flit_output_module1[22]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+22]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[22]));
    MUX21X1 U23(.IN1(head_flit_output_module1[23]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+23]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[23]));
    MUX21X1 U24(.IN1(head_flit_output_module1[24]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+24]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[24]));
    MUX21X1 U25(.IN1(head_flit_output_module1[25]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+25]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[25]));
    MUX21X1 U26(.IN1(head_flit_output_module1[26]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+26]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[26]));
    MUX21X1 U27(.IN1(head_flit_output_module1[27]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+27]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[27]));
    MUX21X1 U28(.IN1(head_flit_output_module1[28]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+28]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[28]));
    MUX21X1 U29(.IN1(head_flit_output_module1[29]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+29]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[29]));
    MUX21X1 U30(.IN1(head_flit_output_module1[30]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+30]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[30]));
    MUX21X1 U31(.IN1(head_flit_output_module1[31]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+31]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[31]));
    MUX21X1 U32(.IN1(head_flit_output_module1[32]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+32]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[32]));
    MUX21X1 U33(.IN1(head_flit_output_module1[33]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+33]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[33]));
    MUX21X1 U34(.IN1(head_flit_output_module1[34]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+34]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[34]));
    MUX21X1 U35(.IN1(head_flit_output_module1[35]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+35]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[35]));
    MUX21X1 U36(.IN1(head_flit_output_module1[36]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+36]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[36]));

    INVX1 U041 ( .A(head_flit_output_module1[32]), .Y(head_flit_output_module1_32_not_output_module1) );
    AND2X1 U1218 ( .IN1(head_flit_output_module1_32_not_output_module1), .IN2(head_flit_output_module1[33]), .Q(and3resu1_output_module1) );
    NOR4X1 U175821 (.IN1(head_flit_output_module1[29]), .IN2(head_flit_output_module1[28]), .IN3(head_flit_output_module1[27]), .IN4(head_flit_output_module1[26]), .Q(nor23resu1_output_module1) );
    NOR4X1 U175831 (.IN1(head_flit_output_module1[25]), .IN2(head_flit_output_module1[24]), .IN3(head_flit_output_module1[23]), .IN4(head_flit_output_module1[22]), .Q(nor23resu2_output_module1) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module1), .IN2(nor23resu2_output_module1), .Q(and4resu1_output_module1) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module1[33]), .IN2(head_flit_output_module1[32]), .Q(nor23resu3_output_module1) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module1), .IN2(and4resu1_output_module1), .Q(and5resu1_output_module1) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module1), .IN2(nor23resu3_output_module1), .Q(or12resu12_output_module1) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[2:1][0]), .IN2(or12resu12_output_module1), .Q(and6resu1_output_module1) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]), .IN2(and6resu1_output_module1), .S(and2resu1_output_module1) ,.Q(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module1[0]),.B(_sv2v_jump_output_module1[1]),.Y(nand1resu_output_module1));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(_sv2v_jump_output_module1_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module1[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module1[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[i_output_module1[1:0] * 4+:4]), .Q(and8resu1_output_module1) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module1[0]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module1[1]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[1]);
    MUX21X1 U3631(.IN1(req_out_output_module1), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(req_out_output_module1);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1[1]), .Q(norfinresu1_output_module1) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module1), .IN2(req_out_output_module1), .Q(and9resu1_output_module1) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module1), .IN2(grant_im_output_module1[(vc_ch_act_out_output_module1 * 4) + i_output_module1[1:0]]), .Q(and10resu1_output_module1) );    

    MUX21X1 U3(.IN1(ext_req_v_o[73:37][3]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+3]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[73:37][4]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+4]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[73:37][5]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+5]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[73:37][6]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+6]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[73:37][7]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+7]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[73:37][8]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+8]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[73:37][9]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+9]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[73:37][10]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+10]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[73:37][11]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+11]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[73:37][12]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+12]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[73:37][13]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+13]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[73:37][14]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+14]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[73:37][15]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+15]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[73:37][16]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+16]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[73:37][17]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+17]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[73:37][18]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+18]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[73:37][19]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+19]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[73:37][20]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+20]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[73:37][21]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+21]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[73:37][22]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+22]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[73:37][23]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+23]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[73:37][24]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+24]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[73:37][25]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+25]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[73:37][26]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+26]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[73:37][27]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+27]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[73:37][28]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+28]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[73:37][29]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+29]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[73:37][30]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+30]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[73:37][31]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+31]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[73:37][32]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+32]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[73:37][33]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+33]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[73:37][34]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+34]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[73:37][35]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+35]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[73:37][36]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+36]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[73:37][0]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[73:37][1]), .IN2(vc_ch_act_out_output_module1[0]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[73:37][2]), .IN2(vc_ch_act_out_output_module1[1]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and11resu1_output_module1) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    
    
 





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter122) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter122[0]), .Y(i_0_not_high_prior_arbiter122) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter122), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter122[0]), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b1), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(_sv2v_jump_high_prior_arbiter122[1]), .QN(nandres_high_prior_arbiter122) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter222[0]), .Y(i_0_not_high_prior_arbiter222) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter222), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter222[0]), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(_sv2v_jump_high_prior_arbiter222[1]), .QN(nandres_high_prior_arbiter222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter22[0]), .B(valid_from_im_output_module2[3:0][0]), .Y(mask_req_rr_arbiter22[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter22[1]), .B(valid_from_im_output_module2[3:0][1]), .Y(mask_req_rr_arbiter22[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter22[0]), .Y(next_mask_rr_arbiter22[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter22[1]), .Y(next_mask_rr_arbiter22[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter22[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter22) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter22[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter22) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter22[0]), .IN2(raw_grant_rr_arbiter22[0]), .S(xnor0res_rr_arbiter22), .Q(grant_im_output_module2[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter22[1]), .IN2(raw_grant_rr_arbiter22[1]), .S(xnor1res_rr_arbiter22), .Q(grant_im_output_module2[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter22[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter22[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter22[1]), .B(1'b0), .Y(firstif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter22), .B(grant_im_output_module2[3:0][i_rr_arbiter22[0]]), .Y(secondif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[1]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter22[0]), .Q(j_rr_arbiter22[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter22), .B(j_rr_arbiter22[0]), .Y(thirdif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[j_rr_arbiter22[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter22), .Q(next_mask_rr_arbiter22[j_rr_arbiter22[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b1), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(_sv2v_jump_rr_rr_arbiter22[1]), .QN(fourthif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter22) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter22) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter22[0]), .IN2(next_mask_rr_arbiter22[0]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter22[1]), .IN2(next_mask_rr_arbiter22[1]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter2222), .IN2(1'sb1), .S(arst_value_rr_arbiter22), .Q(mask_ff_rr_arbiter22[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1221) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1221[0]), .Y(i_0_not_high_prior_arbiter1221) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1221), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1221[0]), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b1), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(_sv2v_jump_high_prior_arbiter1221[1]), .QN(nandres_high_prior_arbiter1221) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22212) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2221[0]), .Y(i_0_not_high_prior_arbiter22212) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22212), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2221[0]), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(_sv2v_jump_high_prior_arbiter2221[1]), .QN(nandres_high_prior_arbiter22212) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter221[0]), .B(valid_from_im_output_module2[7:4][0]), .Y(mask_req_rr_arbiter221[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter221[1]), .B(valid_from_im_output_module2[7:4][1]), .Y(mask_req_rr_arbiter221[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter221[0]), .Y(next_mask_rr_arbiter221[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter221[1]), .Y(next_mask_rr_arbiter221[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter221[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter221) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter221[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter221) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter221[0]), .IN2(raw_grant_rr_arbiter221[0]), .S(xnor0res_rr_arbiter221), .Q(grant_im_output_module2[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter221[1]), .IN2(raw_grant_rr_arbiter221[1]), .S(xnor1res_rr_arbiter221), .Q(grant_im_output_module2[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter221[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter221[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter221[1]), .B(1'b0), .Y(firstif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter221), .B(grant_im_output_module2[7:4][i_rr_arbiter221[0]]), .Y(secondif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[1]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter221[0]), .Q(j_rr_arbiter221[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter221), .B(j_rr_arbiter221[0]), .Y(thirdif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[j_rr_arbiter221[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter221), .Q(next_mask_rr_arbiter221[j_rr_arbiter221[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b1), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(_sv2v_jump_rr_rr_arbiter221[1]), .QN(fourthif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter221) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter221) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter221[0]), .IN2(next_mask_rr_arbiter221[0]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter221[1]), .IN2(next_mask_rr_arbiter221[1]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter222211), .IN2(1'sb1), .S(arst_value_rr_arbiter221), .Q(mask_ff_rr_arbiter221[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1222[0]), .Y(i_0_not_high_prior_arbiter1222) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1222), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1222[0]), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b1), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(_sv2v_jump_high_prior_arbiter1222[1]), .QN(nandres_high_prior_arbiter1222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2222[0]), .Y(i_0_not_high_prior_arbiter2222) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2222), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2222[0]), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(_sv2v_jump_high_prior_arbiter2222[1]), .QN(nandres_high_prior_arbiter2222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter222[0]), .B(valid_from_im_output_module2[11:8][0]), .Y(mask_req_rr_arbiter222[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter222[1]), .B(valid_from_im_output_module2[11:8][1]), .Y(mask_req_rr_arbiter222[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter222[0]), .Y(next_mask_rr_arbiter222[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter222[1]), .Y(next_mask_rr_arbiter222[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter222[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter222) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter222[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter222) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter222[0]), .IN2(raw_grant_rr_arbiter222[0]), .S(xnor0res_rr_arbiter222), .Q(grant_im_output_module2[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter222[1]), .IN2(raw_grant_rr_arbiter222[1]), .S(xnor1res_rr_arbiter222), .Q(grant_im_output_module2[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter222[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter222[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter222[1]), .B(1'b0), .Y(firstif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter222), .B(grant_im_output_module2[11:8][i_rr_arbiter222[0]]), .Y(secondif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[1]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter222[0]), .Q(j_rr_arbiter222[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter222), .B(j_rr_arbiter222[0]), .Y(thirdif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[j_rr_arbiter222[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter222), .Q(next_mask_rr_arbiter222[j_rr_arbiter222[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b1), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(_sv2v_jump_rr_rr_arbiter222[1]), .QN(fourthif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter222) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter222) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter222[0]), .IN2(next_mask_rr_arbiter222[0]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter222[1]), .IN2(next_mask_rr_arbiter222[1]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter222222), .IN2(1'sb1), .S(arst_value_rr_arbiter222), .Q(mask_ff_rr_arbiter222[0]));


    XNOR2X1 U222 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37]), .IN2(vc_channel_output_module2[1]), .QN(xnor1resu1_output_module2) );
    XNOR2X1 U223 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37-1]), .IN2(vc_channel_output_module2[0]), .QN(xnor2resu1_output_module2) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module2), .IN2(xnor2resu1_output_module2), .Q(and1resu1_output_module2) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]), .IN2(1'b1), .S(and1resu1_output_module2), .Q(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .Q(xor1resu1_output_module2) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module2_1[0]), .IN2(_sv2v_jump_output_module2[0]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module2_1[1]), .IN2(_sv2v_jump_output_module2[1]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[vc_channel_output_module2[1:0]*4+in_mod_output_module2[1:0]]), .Q(and2resu1_output_module2) );

    MUX21X1 U3(.IN1(head_flit_output_module2[3]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+3]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[3]));
    MUX21X1 U4(.IN1(head_flit_output_module2[4]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+4]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[4]));
    MUX21X1 U5(.IN1(head_flit_output_module2[5]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+5]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[5]));
    MUX21X1 U6(.IN1(head_flit_output_module2[6]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+6]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[6]));
    MUX21X1 U7(.IN1(head_flit_output_module2[7]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+7]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[7]));
    MUX21X1 U8(.IN1(head_flit_output_module2[8]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+8]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[8]));
    MUX21X1 U9(.IN1(head_flit_output_module2[9]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+9]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[9]));
    MUX21X1 U10(.IN1(head_flit_output_module2[10]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+10]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[10]));
    MUX21X1 U11(.IN1(head_flit_output_module2[11]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+11]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[11]));
    MUX21X1 U12(.IN1(head_flit_output_module2[12]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+12]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[12]));
    MUX21X1 U13(.IN1(head_flit_output_module2[13]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+13]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[13]));
    MUX21X1 U14(.IN1(head_flit_output_module2[14]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+14]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[14]));
    MUX21X1 U15(.IN1(head_flit_output_module2[15]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+15]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[15]));
    MUX21X1 U16(.IN1(head_flit_output_module2[16]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+16]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[16]));
    MUX21X1 U17(.IN1(head_flit_output_module2[17]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+17]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[17]));
    MUX21X1 U18(.IN1(head_flit_output_module2[18]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+18]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[18]));
    MUX21X1 U19(.IN1(head_flit_output_module2[19]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+19]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[19]));
    MUX21X1 U20(.IN1(head_flit_output_module2[20]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+20]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[20]));
    MUX21X1 U21(.IN1(head_flit_output_module2[21]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+21]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[21]));
    MUX21X1 U22(.IN1(head_flit_output_module2[22]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+22]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[22]));
    MUX21X1 U23(.IN1(head_flit_output_module2[23]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+23]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[23]));
    MUX21X1 U24(.IN1(head_flit_output_module2[24]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+24]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[24]));
    MUX21X1 U25(.IN1(head_flit_output_module2[25]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+25]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[25]));
    MUX21X1 U26(.IN1(head_flit_output_module2[26]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+26]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[26]));
    MUX21X1 U27(.IN1(head_flit_output_module2[27]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+27]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[27]));
    MUX21X1 U28(.IN1(head_flit_output_module2[28]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+28]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[28]));
    MUX21X1 U29(.IN1(head_flit_output_module2[29]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+29]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[29]));
    MUX21X1 U30(.IN1(head_flit_output_module2[30]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+30]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[30]));
    MUX21X1 U31(.IN1(head_flit_output_module2[31]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+31]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[31]));
    MUX21X1 U32(.IN1(head_flit_output_module2[32]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+32]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[32]));
    MUX21X1 U33(.IN1(head_flit_output_module2[33]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+33]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[33]));
    MUX21X1 U34(.IN1(head_flit_output_module2[34]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+34]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[34]));
    MUX21X1 U35(.IN1(head_flit_output_module2[35]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+35]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[35]));
    MUX21X1 U36(.IN1(head_flit_output_module2[36]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+36]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[36]));

    INVX1 U041 ( .A(head_flit_output_module2[32]), .Y(head_flit_output_module2_32_not_output_module2) );
    AND2X1 U1218 ( .IN1(head_flit_output_module2_32_not_output_module2), .IN2(head_flit_output_module2[33]), .Q(and3resu1_output_module2) );
    NOR4X1 U175821 (.IN1(head_flit_output_module2[29]), .IN2(head_flit_output_module2[28]), .IN3(head_flit_output_module2[27]), .IN4(head_flit_output_module2[26]), .Q(nor23resu1_output_module2) );
    NOR4X1 U175831 (.IN1(head_flit_output_module2[25]), .IN2(head_flit_output_module2[24]), .IN3(head_flit_output_module2[23]), .IN4(head_flit_output_module2[22]), .Q(nor23resu2_output_module2) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module2), .IN2(nor23resu2_output_module2), .Q(and4resu1_output_module2) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module2[33]), .IN2(head_flit_output_module2[32]), .Q(nor23resu3_output_module2) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module2), .IN2(and4resu1_output_module2), .Q(and5resu1_output_module2) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module2), .IN2(nor23resu3_output_module2), .Q(or12resu12_output_module2) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[3:2][0]), .IN2(or12resu12_output_module2), .Q(and6resu1_output_module2) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]), .IN2(and6resu1_output_module2), .S(and2resu1_output_module2) ,.Q(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module2[0]),.B(_sv2v_jump_output_module2[1]),.Y(nand1resu_output_module2));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(_sv2v_jump_output_module2_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module2[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module2[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[i_output_module2[1:0] * 4+:4]), .Q(and8resu1_output_module2) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module2[0]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module2[1]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[1]);
    MUX21X1 U3631(.IN1(req_out_output_module2), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(req_out_output_module2);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2[1]), .Q(norfinresu1_output_module2) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module2), .IN2(req_out_output_module2), .Q(and9resu1_output_module2) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module2), .IN2(grant_im_output_module2[(vc_ch_act_out_output_module2 * 4) + i_output_module2[1:0]]), .Q(and10resu1_output_module2) );    

    MUX21X1 U3(.IN1(ext_req_v_o[110:74][3]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+3]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[110:74][4]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+4]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[110:74][5]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+5]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[110:74][6]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+6]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[110:74][7]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+7]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[110:74][8]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+8]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[110:74][9]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+9]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[110:74][10]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+10]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[110:74][11]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+11]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[110:74][12]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+12]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[110:74][13]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+13]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[110:74][14]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+14]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[110:74][15]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+15]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[110:74][16]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+16]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[110:74][17]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+17]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[110:74][18]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+18]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[110:74][19]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+19]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[110:74][20]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+20]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[110:74][21]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+21]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[110:74][22]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+22]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[110:74][23]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+23]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[110:74][24]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+24]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[110:74][25]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+25]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[110:74][26]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+26]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[110:74][27]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+27]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[110:74][28]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+28]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[110:74][29]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+29]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[110:74][30]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+30]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[110:74][31]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+31]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[110:74][32]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+32]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[110:74][33]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+33]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[110:74][34]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+34]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[110:74][35]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+35]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[110:74][36]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+36]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[110:74][0]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[110:74][1]), .IN2(vc_ch_act_out_output_module2[0]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[110:74][2]), .IN2(vc_ch_act_out_output_module2[1]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and11resu1_output_module2) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);   










    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter13) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter13[0]), .Y(i_0_not_high_prior_arbiter13) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter13), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter13[0]), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b1), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(_sv2v_jump_high_prior_arbiter13[1]), .QN(nandres_high_prior_arbiter13) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter23) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter23[0]), .Y(i_0_not_high_prior_arbiter23) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter23), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter23[0]), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(_sv2v_jump_high_prior_arbiter23[1]), .QN(nandres_high_prior_arbiter23) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter3[0]), .B(valid_from_im_output_module3[3:0][0]), .Y(mask_req_rr_arbiter3[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter3[1]), .B(valid_from_im_output_module3[3:0][1]), .Y(mask_req_rr_arbiter3[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter3[0]), .Y(next_mask_rr_arbiter3[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter3[1]), .Y(next_mask_rr_arbiter3[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter3[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter3) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter3[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter3) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter3[0]), .IN2(raw_grant_rr_arbiter3[0]), .S(xnor0res_rr_arbiter3), .Q(grant_im_output_module3[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter3[1]), .IN2(raw_grant_rr_arbiter3[1]), .S(xnor1res_rr_arbiter3), .Q(grant_im_output_module3[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter3[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter3[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter3[1]), .B(1'b0), .Y(firstif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter3), .B(grant_im_output_module3[3:0][i_rr_arbiter3[0]]), .Y(secondif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[1]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter3[0]), .Q(j_rr_arbiter3[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter3), .B(j_rr_arbiter3[0]), .Y(thirdif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[j_rr_arbiter3[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter3), .Q(next_mask_rr_arbiter3[j_rr_arbiter3[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b1), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(_sv2v_jump_rr_rr_arbiter3[1]), .QN(fourthif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter3) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter3) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter3[0]), .IN2(next_mask_rr_arbiter3[0]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter3[1]), .IN2(next_mask_rr_arbiter3[1]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter33), .IN2(1'sb1), .S(arst_value_rr_arbiter3), .Q(mask_ff_rr_arbiter3[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter131) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter131[0]), .Y(i_0_not_high_prior_arbiter131) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter131), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter131[0]), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b1), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(_sv2v_jump_high_prior_arbiter131[1]), .QN(nandres_high_prior_arbiter131) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2313) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter231[0]), .Y(i_0_not_high_prior_arbiter2313) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2313), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter231[0]), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(_sv2v_jump_high_prior_arbiter231[1]), .QN(nandres_high_prior_arbiter2313) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter31[0]), .B(valid_from_im_output_module3[7:4][0]), .Y(mask_req_rr_arbiter31[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter31[1]), .B(valid_from_im_output_module3[7:4][1]), .Y(mask_req_rr_arbiter31[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter31[0]), .Y(next_mask_rr_arbiter31[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter31[1]), .Y(next_mask_rr_arbiter31[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter31[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter31) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter31[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter31) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter31[0]), .IN2(raw_grant_rr_arbiter31[0]), .S(xnor0res_rr_arbiter31), .Q(grant_im_output_module3[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter31[1]), .IN2(raw_grant_rr_arbiter31[1]), .S(xnor1res_rr_arbiter31), .Q(grant_im_output_module3[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter31[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter31[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter31[1]), .B(1'b0), .Y(firstif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter31), .B(grant_im_output_module3[7:4][i_rr_arbiter31[0]]), .Y(secondif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[1]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter31[0]), .Q(j_rr_arbiter31[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter31), .B(j_rr_arbiter31[0]), .Y(thirdif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[j_rr_arbiter31[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter31), .Q(next_mask_rr_arbiter31[j_rr_arbiter31[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b1), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(_sv2v_jump_rr_rr_arbiter31[1]), .QN(fourthif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter31) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter31) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter31[0]), .IN2(next_mask_rr_arbiter31[0]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter31[1]), .IN2(next_mask_rr_arbiter31[1]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter3311), .IN2(1'sb1), .S(arst_value_rr_arbiter31), .Q(mask_ff_rr_arbiter31[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter132) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter132[0]), .Y(i_0_not_high_prior_arbiter132) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter132), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter132[0]), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b1), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(_sv2v_jump_high_prior_arbiter132[1]), .QN(nandres_high_prior_arbiter132) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter232) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter232[0]), .Y(i_0_not_high_prior_arbiter232) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter232), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter232[0]), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(_sv2v_jump_high_prior_arbiter232[1]), .QN(nandres_high_prior_arbiter232) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter32[0]), .B(valid_from_im_output_module3[11:8][0]), .Y(mask_req_rr_arbiter32[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter32[1]), .B(valid_from_im_output_module3[11:8][1]), .Y(mask_req_rr_arbiter32[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter32[0]), .Y(next_mask_rr_arbiter32[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter32[1]), .Y(next_mask_rr_arbiter32[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter32[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter32) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter32[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter32) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter32[0]), .IN2(raw_grant_rr_arbiter32[0]), .S(xnor0res_rr_arbiter32), .Q(grant_im_output_module3[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter32[1]), .IN2(raw_grant_rr_arbiter32[1]), .S(xnor1res_rr_arbiter32), .Q(grant_im_output_module3[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter32[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter32[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter32[1]), .B(1'b0), .Y(firstif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter32), .B(grant_im_output_module3[11:8][i_rr_arbiter32[0]]), .Y(secondif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[1]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter32[0]), .Q(j_rr_arbiter32[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter32), .B(j_rr_arbiter32[0]), .Y(thirdif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[j_rr_arbiter32[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter32), .Q(next_mask_rr_arbiter32[j_rr_arbiter32[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b1), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(_sv2v_jump_rr_rr_arbiter32[1]), .QN(fourthif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter32) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter32) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter32[0]), .IN2(next_mask_rr_arbiter32[0]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter32[1]), .IN2(next_mask_rr_arbiter32[1]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter3322), .IN2(1'sb1), .S(arst_value_rr_arbiter32), .Q(mask_ff_rr_arbiter32[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37]), .IN2(vc_channel_output_module3[1]), .QN(xnor1resu1_output_module3) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37-1]), .IN2(vc_channel_output_module3[0]), .QN(xnor2resu1_output_module3) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module3), .IN2(xnor2resu1_output_module3), .Q(and1resu1_output_module3) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]), .IN2(1'b1), .S(and1resu1_output_module3), .Q(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .Q(xor1resu1_output_module3) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module3_1[0]), .IN2(_sv2v_jump_output_module3[0]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module3_1[1]), .IN2(_sv2v_jump_output_module3[1]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[vc_channel_output_module3[1:0]*4+in_mod_output_module3[1:0]]), .Q(and2resu1_output_module3) );

    MUX21X1 U3(.IN1(head_flit_output_module3[3]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+3]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[3]));
    MUX21X1 U4(.IN1(head_flit_output_module3[4]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+4]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[4]));
    MUX21X1 U5(.IN1(head_flit_output_module3[5]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+5]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[5]));
    MUX21X1 U6(.IN1(head_flit_output_module3[6]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+6]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[6]));
    MUX21X1 U7(.IN1(head_flit_output_module3[7]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+7]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[7]));
    MUX21X1 U8(.IN1(head_flit_output_module3[8]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+8]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[8]));
    MUX21X1 U9(.IN1(head_flit_output_module3[9]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+9]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[9]));
    MUX21X1 U10(.IN1(head_flit_output_module3[10]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+10]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[10]));
    MUX21X1 U11(.IN1(head_flit_output_module3[11]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+11]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[11]));
    MUX21X1 U12(.IN1(head_flit_output_module3[12]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+12]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[12]));
    MUX21X1 U13(.IN1(head_flit_output_module3[13]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+13]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[13]));
    MUX21X1 U14(.IN1(head_flit_output_module3[14]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+14]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[14]));
    MUX21X1 U15(.IN1(head_flit_output_module3[15]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+15]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[15]));
    MUX21X1 U16(.IN1(head_flit_output_module3[16]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+16]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[16]));
    MUX21X1 U17(.IN1(head_flit_output_module3[17]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+17]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[17]));
    MUX21X1 U18(.IN1(head_flit_output_module3[18]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+18]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[18]));
    MUX21X1 U19(.IN1(head_flit_output_module3[19]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+19]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[19]));
    MUX21X1 U20(.IN1(head_flit_output_module3[20]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+20]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[20]));
    MUX21X1 U21(.IN1(head_flit_output_module3[21]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+21]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[21]));
    MUX21X1 U22(.IN1(head_flit_output_module3[22]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+22]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[22]));
    MUX21X1 U23(.IN1(head_flit_output_module3[23]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+23]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[23]));
    MUX21X1 U24(.IN1(head_flit_output_module3[24]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+24]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[24]));
    MUX21X1 U25(.IN1(head_flit_output_module3[25]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+25]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[25]));
    MUX21X1 U26(.IN1(head_flit_output_module3[26]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+26]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[26]));
    MUX21X1 U27(.IN1(head_flit_output_module3[27]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+27]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[27]));
    MUX21X1 U28(.IN1(head_flit_output_module3[28]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+28]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[28]));
    MUX21X1 U29(.IN1(head_flit_output_module3[29]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+29]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[29]));
    MUX21X1 U30(.IN1(head_flit_output_module3[30]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+30]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[30]));
    MUX21X1 U31(.IN1(head_flit_output_module3[31]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+31]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[31]));
    MUX21X1 U32(.IN1(head_flit_output_module3[32]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+32]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[32]));
    MUX21X1 U33(.IN1(head_flit_output_module3[33]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+33]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[33]));
    MUX21X1 U34(.IN1(head_flit_output_module3[34]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+34]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[34]));
    MUX21X1 U35(.IN1(head_flit_output_module3[35]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+35]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[35]));
    MUX21X1 U36(.IN1(head_flit_output_module3[36]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+36]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[36]));

    INVX1 U041 ( .A(head_flit_output_module3[32]), .Y(head_flit_output_module3_32_not_output_module3) );
    AND2X1 U1218 ( .IN1(head_flit_output_module3_32_not_output_module3), .IN2(head_flit_output_module3[33]), .Q(and3resu1_output_module3) );
    NOR4X1 U175821 (.IN1(head_flit_output_module3[29]), .IN2(head_flit_output_module3[28]), .IN3(head_flit_output_module3[27]), .IN4(head_flit_output_module3[26]), .Q(nor23resu1_output_module3) );
    NOR4X1 U175831 (.IN1(head_flit_output_module3[25]), .IN2(head_flit_output_module3[24]), .IN3(head_flit_output_module3[23]), .IN4(head_flit_output_module3[22]), .Q(nor23resu2_output_module3) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module3), .IN2(nor23resu2_output_module3), .Q(and4resu1_output_module3) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module3[33]), .IN2(head_flit_output_module3[32]), .Q(nor23resu3_output_module3) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module3), .IN2(and4resu1_output_module3), .Q(and5resu1_output_module3) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module3), .IN2(nor23resu3_output_module3), .Q(or12resu12_output_module3) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[4:3][0]), .IN2(or12resu12_output_module3), .Q(and6resu1_output_module3) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]), .IN2(and6resu1_output_module3), .S(and2resu1_output_module3) ,.Q(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module3[0]),.B(_sv2v_jump_output_module3[1]),.Y(nand1resu_output_module3));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(_sv2v_jump_output_module3_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module3[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module3[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[i_output_module3[1:0] * 4+:4]), .Q(and8resu1_output_module3) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module3[0]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module3[1]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[1]);
    MUX21X1 U3631(.IN1(req_out_output_module3), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(req_out_output_module3);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3[1]), .Q(norfinresu1_output_module3) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module3), .IN2(req_out_output_module3), .Q(and9resu1_output_module3) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module3), .IN2(grant_im_output_module3[(vc_ch_act_out_output_module3 * 4) + i_output_module3[1:0]]), .Q(and10resu1_output_module3) );    

    MUX21X1 U3(.IN1(ext_req_v_o[147:111][3]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+3]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[147:111][4]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+4]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[147:111][5]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+5]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[147:111][6]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+6]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[147:111][7]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+7]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[147:111][8]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+8]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[147:111][9]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+9]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[147:111][10]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+10]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[147:111][11]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+11]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[147:111][12]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+12]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[147:111][13]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+13]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[147:111][14]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+14]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[147:111][15]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+15]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[147:111][16]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+16]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[147:111][17]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+17]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[147:111][18]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+18]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[147:111][19]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+19]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[147:111][20]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+20]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[147:111][21]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+21]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[147:111][22]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+22]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[147:111][23]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+23]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[147:111][24]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+24]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[147:111][25]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+25]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[147:111][26]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+26]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[147:111][27]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+27]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[147:111][28]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+28]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[147:111][29]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+29]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[147:111][30]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+30]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[147:111][31]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+31]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[147:111][32]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+32]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[147:111][33]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+33]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[147:111][34]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+34]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[147:111][35]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+35]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[147:111][36]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+36]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[147:111][0]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[147:111][1]), .IN2(vc_ch_act_out_output_module3[0]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[147:111][2]), .IN2(vc_ch_act_out_output_module3[1]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and11resu1_output_module3) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    







    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter14) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter14[0]), .Y(i_0_not_high_prior_arbiter14) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter14), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter14[0]), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b1), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(_sv2v_jump_high_prior_arbiter14[1]), .QN(nandres_high_prior_arbiter14) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter24) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter24[0]), .Y(i_0_not_high_prior_arbiter24) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter24), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter24[0]), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(_sv2v_jump_high_prior_arbiter24[1]), .QN(nandres_high_prior_arbiter24) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter4[0]), .B(valid_from_im_output_module4[3:0][0]), .Y(mask_req_rr_arbiter4[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter4[1]), .B(valid_from_im_output_module4[3:0][1]), .Y(mask_req_rr_arbiter4[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter4[0]), .Y(next_mask_rr_arbiter4[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter4[1]), .Y(next_mask_rr_arbiter4[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter4[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter4) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter4[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter4) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter4[0]), .IN2(raw_grant_rr_arbiter4[0]), .S(xnor0res_rr_arbiter4), .Q(grant_im_output_module4[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter4[1]), .IN2(raw_grant_rr_arbiter4[1]), .S(xnor1res_rr_arbiter4), .Q(grant_im_output_module4[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter4[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter4[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter4[1]), .B(1'b0), .Y(firstif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter4), .B(grant_im_output_module4[3:0][i_rr_arbiter4[0]]), .Y(secondif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[1]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter4[0]), .Q(j_rr_arbiter4[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter4), .B(j_rr_arbiter4[0]), .Y(thirdif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[j_rr_arbiter4[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter4), .Q(next_mask_rr_arbiter4[j_rr_arbiter4[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b1), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(_sv2v_jump_rr_rr_arbiter4[1]), .QN(fourthif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter4) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter4) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter4[0]), .IN2(next_mask_rr_arbiter4[0]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter4[1]), .IN2(next_mask_rr_arbiter4[1]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter44), .IN2(1'sb1), .S(arst_value_rr_arbiter4), .Q(mask_ff_rr_arbiter4[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter141) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter141[0]), .Y(i_0_not_high_prior_arbiter141) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter141), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter141[0]), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b1), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(_sv2v_jump_high_prior_arbiter141[1]), .QN(nandres_high_prior_arbiter141) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2414) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter241[0]), .Y(i_0_not_high_prior_arbiter2414) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2414), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter241[0]), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(_sv2v_jump_high_prior_arbiter241[1]), .QN(nandres_high_prior_arbiter2414) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter41[0]), .B(valid_from_im_output_module4[7:4][0]), .Y(mask_req_rr_arbiter41[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter41[1]), .B(valid_from_im_output_module4[7:4][1]), .Y(mask_req_rr_arbiter41[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter41[0]), .Y(next_mask_rr_arbiter41[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter41[1]), .Y(next_mask_rr_arbiter41[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter41[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter41) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter41[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter41) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter41[0]), .IN2(raw_grant_rr_arbiter41[0]), .S(xnor0res_rr_arbiter41), .Q(grant_im_output_module4[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter41[1]), .IN2(raw_grant_rr_arbiter41[1]), .S(xnor1res_rr_arbiter41), .Q(grant_im_output_module4[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter41[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter41[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter41[1]), .B(1'b0), .Y(firstif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter41), .B(grant_im_output_module4[7:4][i_rr_arbiter41[0]]), .Y(secondif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[1]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter41[0]), .Q(j_rr_arbiter41[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter41), .B(j_rr_arbiter41[0]), .Y(thirdif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[j_rr_arbiter41[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter41), .Q(next_mask_rr_arbiter41[j_rr_arbiter41[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b1), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(_sv2v_jump_rr_rr_arbiter41[1]), .QN(fourthif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter41) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter41) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter41[0]), .IN2(next_mask_rr_arbiter41[0]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter41[1]), .IN2(next_mask_rr_arbiter41[1]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter4411), .IN2(1'sb1), .S(arst_value_rr_arbiter41), .Q(mask_ff_rr_arbiter41[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter142) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter142[0]), .Y(i_0_not_high_prior_arbiter142) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter142), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter142[0]), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b1), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(_sv2v_jump_high_prior_arbiter142[1]), .QN(nandres_high_prior_arbiter142) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter242) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter242[0]), .Y(i_0_not_high_prior_arbiter242) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter242), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter242[0]), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(_sv2v_jump_high_prior_arbiter242[1]), .QN(nandres_high_prior_arbiter242) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter42[0]), .B(valid_from_im_output_module4[11:8][0]), .Y(mask_req_rr_arbiter42[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter42[1]), .B(valid_from_im_output_module4[11:8][1]), .Y(mask_req_rr_arbiter42[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter42[0]), .Y(next_mask_rr_arbiter42[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter42[1]), .Y(next_mask_rr_arbiter42[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter42[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter42) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter42[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter42) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter42[0]), .IN2(raw_grant_rr_arbiter42[0]), .S(xnor0res_rr_arbiter42), .Q(grant_im_output_module4[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter42[1]), .IN2(raw_grant_rr_arbiter42[1]), .S(xnor1res_rr_arbiter42), .Q(grant_im_output_module4[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter42[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter42[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter42[1]), .B(1'b0), .Y(firstif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter42), .B(grant_im_output_module4[11:8][i_rr_arbiter42[0]]), .Y(secondif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[1]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter42[0]), .Q(j_rr_arbiter42[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter42), .B(j_rr_arbiter42[0]), .Y(thirdif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[j_rr_arbiter42[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter42), .Q(next_mask_rr_arbiter42[j_rr_arbiter42[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b1), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(_sv2v_jump_rr_rr_arbiter42[1]), .QN(fourthif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter42) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter42) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter42[0]), .IN2(next_mask_rr_arbiter42[0]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter42[1]), .IN2(next_mask_rr_arbiter42[1]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter4422), .IN2(1'sb1), .S(arst_value_rr_arbiter42), .Q(mask_ff_rr_arbiter42[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37]), .IN2(vc_channel_output_module4[1]), .QN(xnor1resu1_output_module4) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37-1]), .IN2(vc_channel_output_module4[0]), .QN(xnor2resu1_output_module4) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module4), .IN2(xnor2resu1_output_module4), .Q(and1resu1_output_module4) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]), .IN2(1'b1), .S(and1resu1_output_module4), .Q(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .Q(xor1resu1_output_module4) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module4_1[0]), .IN2(_sv2v_jump_output_module4[0]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module4_1[1]), .IN2(_sv2v_jump_output_module4[1]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[vc_channel_output_module4[1:0]*4+in_mod_output_module4[1:0]]), .Q(and2resu1_output_module4) );

    MUX21X1 U3(.IN1(head_flit_output_module4[3]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+3]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[3]));
    MUX21X1 U4(.IN1(head_flit_output_module4[4]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+4]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[4]));
    MUX21X1 U5(.IN1(head_flit_output_module4[5]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+5]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[5]));
    MUX21X1 U6(.IN1(head_flit_output_module4[6]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+6]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[6]));
    MUX21X1 U7(.IN1(head_flit_output_module4[7]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+7]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[7]));
    MUX21X1 U8(.IN1(head_flit_output_module4[8]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+8]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[8]));
    MUX21X1 U9(.IN1(head_flit_output_module4[9]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+9]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[9]));
    MUX21X1 U10(.IN1(head_flit_output_module4[10]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+10]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[10]));
    MUX21X1 U11(.IN1(head_flit_output_module4[11]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+11]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[11]));
    MUX21X1 U12(.IN1(head_flit_output_module4[12]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+12]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[12]));
    MUX21X1 U13(.IN1(head_flit_output_module4[13]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+13]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[13]));
    MUX21X1 U14(.IN1(head_flit_output_module4[14]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+14]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[14]));
    MUX21X1 U15(.IN1(head_flit_output_module4[15]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+15]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[15]));
    MUX21X1 U16(.IN1(head_flit_output_module4[16]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+16]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[16]));
    MUX21X1 U17(.IN1(head_flit_output_module4[17]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+17]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[17]));
    MUX21X1 U18(.IN1(head_flit_output_module4[18]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+18]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[18]));
    MUX21X1 U19(.IN1(head_flit_output_module4[19]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+19]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[19]));
    MUX21X1 U20(.IN1(head_flit_output_module4[20]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+20]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[20]));
    MUX21X1 U21(.IN1(head_flit_output_module4[21]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+21]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[21]));
    MUX21X1 U22(.IN1(head_flit_output_module4[22]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+22]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[22]));
    MUX21X1 U23(.IN1(head_flit_output_module4[23]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+23]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[23]));
    MUX21X1 U24(.IN1(head_flit_output_module4[24]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+24]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[24]));
    MUX21X1 U25(.IN1(head_flit_output_module4[25]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+25]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[25]));
    MUX21X1 U26(.IN1(head_flit_output_module4[26]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+26]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[26]));
    MUX21X1 U27(.IN1(head_flit_output_module4[27]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+27]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[27]));
    MUX21X1 U28(.IN1(head_flit_output_module4[28]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+28]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[28]));
    MUX21X1 U29(.IN1(head_flit_output_module4[29]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+29]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[29]));
    MUX21X1 U30(.IN1(head_flit_output_module4[30]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+30]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[30]));
    MUX21X1 U31(.IN1(head_flit_output_module4[31]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+31]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[31]));
    MUX21X1 U32(.IN1(head_flit_output_module4[32]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+32]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[32]));
    MUX21X1 U33(.IN1(head_flit_output_module4[33]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+33]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[33]));
    MUX21X1 U34(.IN1(head_flit_output_module4[34]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+34]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[34]));
    MUX21X1 U35(.IN1(head_flit_output_module4[35]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+35]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[35]));
    MUX21X1 U36(.IN1(head_flit_output_module4[36]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+36]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[36]));

    INVX1 U041 ( .A(head_flit_output_module4[32]), .Y(head_flit_output_module4_32_not_output_module4) );
    AND2X1 U1218 ( .IN1(head_flit_output_module4_32_not_output_module4), .IN2(head_flit_output_module4[33]), .Q(and3resu1_output_module4) );
    NOR4X1 U175821 (.IN1(head_flit_output_module4[29]), .IN2(head_flit_output_module4[28]), .IN3(head_flit_output_module4[27]), .IN4(head_flit_output_module4[26]), .Q(nor23resu1_output_module4) );
    NOR4X1 U175831 (.IN1(head_flit_output_module4[25]), .IN2(head_flit_output_module4[24]), .IN3(head_flit_output_module4[23]), .IN4(head_flit_output_module4[22]), .Q(nor23resu2_output_module4) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module4), .IN2(nor23resu2_output_module4), .Q(and4resu1_output_module4) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module4[33]), .IN2(head_flit_output_module4[32]), .Q(nor23resu3_output_module4) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module4), .IN2(and4resu1_output_module4), .Q(and5resu1_output_module4) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module4), .IN2(nor23resu3_output_module4), .Q(or12resu12_output_module4) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[5:4][0]), .IN2(or12resu12_output_module4), .Q(and6resu1_output_module4) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]), .IN2(and6resu1_output_module4), .S(and2resu1_output_module4) ,.Q(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module4[0]),.B(_sv2v_jump_output_module4[1]),.Y(nand1resu_output_module4));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(_sv2v_jump_output_module4_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module4[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module4[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[i_output_module4[1:0] * 4+:4]), .Q(and8resu1_output_module4) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module4[0]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module4[1]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[1]);
    MUX21X1 U3631(.IN1(req_out_output_module4), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(req_out_output_module4);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4[1]), .Q(norfinresu1_output_module4) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module4), .IN2(req_out_output_module4), .Q(and9resu1_output_module4) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module4), .IN2(grant_im_output_module4[(vc_ch_act_out_output_module4 * 4) + i_output_module4[1:0]]), .Q(and10resu1_output_module4) );    

    MUX21X1 U3(.IN1(ext_req_v_o[184:148][3]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+3]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[184:148][4]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+4]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[184:148][5]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+5]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[184:148][6]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+6]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[184:148][7]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+7]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[184:148][8]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+8]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[184:148][9]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+9]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[184:148][10]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+10]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[184:148][11]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+11]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[184:148][12]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+12]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[184:148][13]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+13]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[184:148][14]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+14]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[184:148][15]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+15]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[184:148][16]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+16]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[184:148][17]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+17]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[184:148][18]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+18]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[184:148][19]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+19]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[184:148][20]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+20]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[184:148][21]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+21]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[184:148][22]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+22]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[184:148][23]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+23]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[184:148][24]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+24]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[184:148][25]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+25]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[184:148][26]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+26]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[184:148][27]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+27]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[184:148][28]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+28]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[184:148][29]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+29]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[184:148][30]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+30]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[184:148][31]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+31]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[184:148][32]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+32]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[184:148][33]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+33]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[184:148][34]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+34]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[184:148][35]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+35]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[184:148][36]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+36]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[184:148][0]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[184:148][1]), .IN2(vc_ch_act_out_output_module4[0]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[184:148][2]), .IN2(vc_ch_act_out_output_module4[1]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and11resu1_output_module4) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    



//router body
	BUFX1 U001 ( .A(north_recv_req), .Y(ext_req_v_i[0]) );
	BUFX1 U002 ( .A(north_recv_resp), .Y(ext_resp_v_o[0]) );
	BUFX1 U003 ( .A(xt_req_v_i[37]), .Y(south_recv_req) );
	BUFX1 U004 ( .A(south_recv_resp), .Y(ext_resp_v_o[1]) );
	BUFX1 U005 ( .A(ext_req_v_i[74]), .Y(west_recv_req) );
	BUFX1 U006 ( .A(west_recv_resp), .Y(ext_resp_v_o[2]) );
	BUFX1 U007 ( .A(ext_req_v_i[111]), .Y(east_recv_req) );
	BUFX1 U008 ( .A(east_recv_resp), .Y(ext_resp_v_o[3]) );
	BUFX1 U009 ( .A(north_send_req), .Y(ext_req_v_o[0]) );
	BUFX1 U010 ( .A(ext_resp_v_i[0]), .Y(north_send_resp) );
	BUFX1 U011 ( .A(south_send_req), .Y(ext_req_v_o[37]) );
	BUFX1 U012 ( .A(ext_resp_v_i[1]), .Y(south_send_resp) );
	BUFX1 U013 ( .A(west_send_req), .Y(ext_req_v_o[74]) );
	BUFX1 U014 ( .A(ext_resp_v_i[2]), .Y(west_send_resp) );
	BUFX1 U015 ( .A(east_send_req), .Y(ext_req_v_o[111]) );
	BUFX1 U016 ( .A(ext_resp_v_i[3]), .Y(east_send_resp) );
	BUFX1 U017 ( .A(local_recv_resp), .Y(ext_resp_v_o[4]) );
	BUFX1 U018 ( .A(ext_req_v_i[148]), .Y(local_recv_req) );
	BUFX1 U019 ( .A(local_send_req), .Y(ext_req_v_o[148]) );
	BUFX1 U020 ( .A(ext_resp_v_i[4]), .Y(local_send_resp) );


	MUX21X1 U0(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[24]) ,.Q(int_map_req_v[0]));
	MUX21X1 U1(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[24]) ,.Q(int_map_req_v[1]));
	MUX21X1 U2(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[24]) ,.Q(int_map_req_v[2]));
	MUX21X1 U3(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[24]) ,.Q(int_map_req_v[3]));
	MUX21X1 U4(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[24]) ,.Q(int_map_req_v[4]));
	MUX21X1 U5(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[24]) ,.Q(int_map_req_v[5]));
	MUX21X1 U6(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[24]) ,.Q(int_map_req_v[6]));
	MUX21X1 U7(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[24]) ,.Q(int_map_req_v[7]));
	MUX21X1 U8(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[24]) ,.Q(int_map_req_v[8]));
	MUX21X1 U9(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[24]) ,.Q(int_map_req_v[9]));
	MUX21X1 U10(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[24]) ,.Q(int_map_req_v[10]));
	MUX21X1 U11(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[24]) ,.Q(int_map_req_v[11]));
	MUX21X1 U12(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[24]) ,.Q(int_map_req_v[12]));
	MUX21X1 U13(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[24]) ,.Q(int_map_req_v[13]));
	MUX21X1 U14(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[24]) ,.Q(int_map_req_v[14]));
	MUX21X1 U15(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[24]) ,.Q(int_map_req_v[15]));
	MUX21X1 U16(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[24]) ,.Q(int_map_req_v[16]));
	MUX21X1 U17(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[24]) ,.Q(int_map_req_v[17]));
	MUX21X1 U18(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[24]) ,.Q(int_map_req_v[18]));
	MUX21X1 U19(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[24]) ,.Q(int_map_req_v[19]));
	MUX21X1 U20(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[24]) ,.Q(int_map_req_v[20]));
	MUX21X1 U21(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[24]) ,.Q(int_map_req_v[21]));
	MUX21X1 U22(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[24]) ,.Q(int_map_req_v[22]));
	MUX21X1 U23(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[24]) ,.Q(int_map_req_v[23]));
	MUX21X1 U24(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[24]) ,.Q(int_map_req_v[24]));
	MUX21X1 U25(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[24]) ,.Q(int_map_req_v[25]));
	MUX21X1 U26(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[24]) ,.Q(int_map_req_v[26]));
	MUX21X1 U27(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[24]) ,.Q(int_map_req_v[27]));
	MUX21X1 U28(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[24]) ,.Q(int_map_req_v[28]));
	MUX21X1 U29(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[24]) ,.Q(int_map_req_v[29]));
	MUX21X1 U30(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[24]) ,.Q(int_map_req_v[30]));
	MUX21X1 U31(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[24]) ,.Q(int_map_req_v[31]));
	MUX21X1 U32(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[24]) ,.Q(int_map_req_v[32]));
	MUX21X1 U33(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[24]) ,.Q(int_map_req_v[33]));
	MUX21X1 U34(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[24]) ,.Q(int_map_req_v[34]));
	MUX21X1 U35(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[24]) ,.Q(int_map_req_v[35]));
	MUX21X1 U36(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[24]) ,.Q(int_map_req_v[36]));
	MUX21X1 U37(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[19]) ,.Q(int_map_req_v[37]));
	MUX21X1 U38(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[19]) ,.Q(int_map_req_v[38]));
	MUX21X1 U39(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[19]) ,.Q(int_map_req_v[39]));
	MUX21X1 U40(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[19]) ,.Q(int_map_req_v[40]));
	MUX21X1 U41(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[19]) ,.Q(int_map_req_v[41]));
	MUX21X1 U42(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[19]) ,.Q(int_map_req_v[42]));
	MUX21X1 U43(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[19]) ,.Q(int_map_req_v[43]));
	MUX21X1 U44(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[19]) ,.Q(int_map_req_v[44]));
	MUX21X1 U45(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[19]) ,.Q(int_map_req_v[45]));
	MUX21X1 U46(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[19]) ,.Q(int_map_req_v[46]));
	MUX21X1 U47(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[19]) ,.Q(int_map_req_v[47]));
	MUX21X1 U48(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[19]) ,.Q(int_map_req_v[48]));
	MUX21X1 U49(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[19]) ,.Q(int_map_req_v[49]));
	MUX21X1 U50(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[19]) ,.Q(int_map_req_v[50]));
	MUX21X1 U51(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[19]) ,.Q(int_map_req_v[51]));
	MUX21X1 U52(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[19]) ,.Q(int_map_req_v[52]));
	MUX21X1 U53(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[19]) ,.Q(int_map_req_v[53]));
	MUX21X1 U54(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[19]) ,.Q(int_map_req_v[54]));
	MUX21X1 U55(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[19]) ,.Q(int_map_req_v[55]));
	MUX21X1 U56(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[19]) ,.Q(int_map_req_v[56]));
	MUX21X1 U57(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[19]) ,.Q(int_map_req_v[57]));
	MUX21X1 U58(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[19]) ,.Q(int_map_req_v[58]));
	MUX21X1 U59(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[19]) ,.Q(int_map_req_v[59]));
	MUX21X1 U60(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[19]) ,.Q(int_map_req_v[60]));
	MUX21X1 U61(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[19]) ,.Q(int_map_req_v[61]));
	MUX21X1 U62(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[19]) ,.Q(int_map_req_v[62]));
	MUX21X1 U63(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[19]) ,.Q(int_map_req_v[63]));
	MUX21X1 U64(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[19]) ,.Q(int_map_req_v[64]));
	MUX21X1 U65(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[19]) ,.Q(int_map_req_v[65]));
	MUX21X1 U66(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[19]) ,.Q(int_map_req_v[66]));
	MUX21X1 U67(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[19]) ,.Q(int_map_req_v[67]));
	MUX21X1 U68(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[19]) ,.Q(int_map_req_v[68]));
	MUX21X1 U69(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[19]) ,.Q(int_map_req_v[69]));
	MUX21X1 U70(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[19]) ,.Q(int_map_req_v[70]));
	MUX21X1 U71(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[19]) ,.Q(int_map_req_v[71]));
	MUX21X1 U72(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[19]) ,.Q(int_map_req_v[72]));
	MUX21X1 U73(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[19]) ,.Q(int_map_req_v[73]));
	MUX21X1 U74(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[14]) ,.Q(int_map_req_v[74]));
	MUX21X1 U75(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[14]) ,.Q(int_map_req_v[75]));
	MUX21X1 U76(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[14]) ,.Q(int_map_req_v[76]));
	MUX21X1 U77(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[14]) ,.Q(int_map_req_v[77]));
	MUX21X1 U78(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[14]) ,.Q(int_map_req_v[78]));
	MUX21X1 U79(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[14]) ,.Q(int_map_req_v[79]));
	MUX21X1 U80(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[14]) ,.Q(int_map_req_v[80]));
	MUX21X1 U81(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[14]) ,.Q(int_map_req_v[81]));
	MUX21X1 U82(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[14]) ,.Q(int_map_req_v[82]));
	MUX21X1 U83(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[14]) ,.Q(int_map_req_v[83]));
	MUX21X1 U84(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[14]) ,.Q(int_map_req_v[84]));
	MUX21X1 U85(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[14]) ,.Q(int_map_req_v[85]));
	MUX21X1 U86(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[14]) ,.Q(int_map_req_v[86]));
	MUX21X1 U87(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[14]) ,.Q(int_map_req_v[87]));
	MUX21X1 U88(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[14]) ,.Q(int_map_req_v[88]));
	MUX21X1 U89(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[14]) ,.Q(int_map_req_v[89]));
	MUX21X1 U90(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[14]) ,.Q(int_map_req_v[90]));
	MUX21X1 U91(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[14]) ,.Q(int_map_req_v[91]));
	MUX21X1 U92(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[14]) ,.Q(int_map_req_v[92]));
	MUX21X1 U93(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[14]) ,.Q(int_map_req_v[93]));
	MUX21X1 U94(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[14]) ,.Q(int_map_req_v[94]));
	MUX21X1 U95(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[14]) ,.Q(int_map_req_v[95]));
	MUX21X1 U96(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[14]) ,.Q(int_map_req_v[96]));
	MUX21X1 U97(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[14]) ,.Q(int_map_req_v[97]));
	MUX21X1 U98(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[14]) ,.Q(int_map_req_v[98]));
	MUX21X1 U99(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[14]) ,.Q(int_map_req_v[99]));
	MUX21X1 U100(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[14]) ,.Q(int_map_req_v[100]));
	MUX21X1 U101(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[14]) ,.Q(int_map_req_v[101]));
	MUX21X1 U102(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[14]) ,.Q(int_map_req_v[102]));
	MUX21X1 U103(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[14]) ,.Q(int_map_req_v[103]));
	MUX21X1 U104(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[14]) ,.Q(int_map_req_v[104]));
	MUX21X1 U105(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[14]) ,.Q(int_map_req_v[105]));
	MUX21X1 U106(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[14]) ,.Q(int_map_req_v[106]));
	MUX21X1 U107(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[14]) ,.Q(int_map_req_v[107]));
	MUX21X1 U108(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[14]) ,.Q(int_map_req_v[108]));
	MUX21X1 U109(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[14]) ,.Q(int_map_req_v[109]));
	MUX21X1 U110(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[14]) ,.Q(int_map_req_v[110]));
	MUX21X1 U111(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[9]) ,.Q(int_map_req_v[111]));
	MUX21X1 U112(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[9]) ,.Q(int_map_req_v[112]));
	MUX21X1 U113(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[9]) ,.Q(int_map_req_v[113]));
	MUX21X1 U114(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[9]) ,.Q(int_map_req_v[114]));
	MUX21X1 U115(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[9]) ,.Q(int_map_req_v[115]));
	MUX21X1 U116(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[9]) ,.Q(int_map_req_v[116]));
	MUX21X1 U117(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[9]) ,.Q(int_map_req_v[117]));
	MUX21X1 U118(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[9]) ,.Q(int_map_req_v[118]));
	MUX21X1 U119(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[9]) ,.Q(int_map_req_v[119]));
	MUX21X1 U120(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[9]) ,.Q(int_map_req_v[120]));
	MUX21X1 U121(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[9]) ,.Q(int_map_req_v[121]));
	MUX21X1 U122(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[9]) ,.Q(int_map_req_v[122]));
	MUX21X1 U123(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[9]) ,.Q(int_map_req_v[123]));
	MUX21X1 U124(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[9]) ,.Q(int_map_req_v[124]));
	MUX21X1 U125(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[9]) ,.Q(int_map_req_v[125]));
	MUX21X1 U126(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[9]) ,.Q(int_map_req_v[126]));
	MUX21X1 U127(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[9]) ,.Q(int_map_req_v[127]));
	MUX21X1 U128(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[9]) ,.Q(int_map_req_v[128]));
	MUX21X1 U129(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[9]) ,.Q(int_map_req_v[129]));
	MUX21X1 U130(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[9]) ,.Q(int_map_req_v[130]));
	MUX21X1 U131(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[9]) ,.Q(int_map_req_v[131]));
	MUX21X1 U132(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[9]) ,.Q(int_map_req_v[132]));
	MUX21X1 U133(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[9]) ,.Q(int_map_req_v[133]));
	MUX21X1 U134(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[9]) ,.Q(int_map_req_v[134]));
	MUX21X1 U135(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[9]) ,.Q(int_map_req_v[135]));
	MUX21X1 U136(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[9]) ,.Q(int_map_req_v[136]));
	MUX21X1 U137(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[9]) ,.Q(int_map_req_v[137]));
	MUX21X1 U138(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[9]) ,.Q(int_map_req_v[138]));
	MUX21X1 U139(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[9]) ,.Q(int_map_req_v[139]));
	MUX21X1 U140(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[9]) ,.Q(int_map_req_v[140]));
	MUX21X1 U141(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[9]) ,.Q(int_map_req_v[141]));
	MUX21X1 U142(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[9]) ,.Q(int_map_req_v[142]));
	MUX21X1 U143(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[9]) ,.Q(int_map_req_v[143]));
	MUX21X1 U144(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[9]) ,.Q(int_map_req_v[144]));
	MUX21X1 U145(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[9]) ,.Q(int_map_req_v[145]));
	MUX21X1 U146(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[9]) ,.Q(int_map_req_v[146]));
	MUX21X1 U147(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[9]) ,.Q(int_map_req_v[147]));
	MUX21X1 U01(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[3]), .S(int_route_v[9]) ,.Q(int_resp_v[1]));
	MUX21X1 U02(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[4]), .S(int_route_v[9]) ,.Q(int_resp_v[2]));
	MUX21X1 U03(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[2]), .S(int_route_v[14]) ,.Q(int_resp_v[2]));
	MUX21X1 U04(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[3]), .S(int_route_v[14]) ,.Q(int_resp_v[3]));
	MUX21X1 U05(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[1]), .S(int_route_v[19]) ,.Q(int_resp_v[3]));
	MUX21X1 U06(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[2]), .S(int_route_v[19]) ,.Q(int_resp_v[4]));
	MUX21X1 U07(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[0]), .S(int_route_v[24]) ,.Q(int_resp_v[4]));
	MUX21X1 U08(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[1]), .S(int_route_v[24]) ,.Q(int_resp_v[5]));


	MUX21X1 U148(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[3]) ,.Q(int_map_req_v[148]));
	MUX21X1 U149(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[3]) ,.Q(int_map_req_v[149]));
	MUX21X1 U150(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[3]) ,.Q(int_map_req_v[150]));
	MUX21X1 U151(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[3]) ,.Q(int_map_req_v[151]));
	MUX21X1 U152(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[3]) ,.Q(int_map_req_v[152]));
	MUX21X1 U153(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[3]) ,.Q(int_map_req_v[153]));
	MUX21X1 U154(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[3]) ,.Q(int_map_req_v[154]));
	MUX21X1 U155(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[3]) ,.Q(int_map_req_v[155]));
	MUX21X1 U156(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[3]) ,.Q(int_map_req_v[156]));
	MUX21X1 U157(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[3]) ,.Q(int_map_req_v[157]));
	MUX21X1 U158(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[3]) ,.Q(int_map_req_v[158]));
	MUX21X1 U159(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[3]) ,.Q(int_map_req_v[159]));
	MUX21X1 U160(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[3]) ,.Q(int_map_req_v[160]));
	MUX21X1 U161(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[3]) ,.Q(int_map_req_v[161]));
	MUX21X1 U162(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[3]) ,.Q(int_map_req_v[162]));
	MUX21X1 U163(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[3]) ,.Q(int_map_req_v[163]));
	MUX21X1 U164(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[3]) ,.Q(int_map_req_v[164]));
	MUX21X1 U165(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[3]) ,.Q(int_map_req_v[165]));
	MUX21X1 U166(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[3]) ,.Q(int_map_req_v[166]));
	MUX21X1 U167(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[3]) ,.Q(int_map_req_v[167]));
	MUX21X1 U168(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[3]) ,.Q(int_map_req_v[168]));
	MUX21X1 U169(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[3]) ,.Q(int_map_req_v[169]));
	MUX21X1 U170(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[3]) ,.Q(int_map_req_v[170]));
	MUX21X1 U171(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[3]) ,.Q(int_map_req_v[171]));
	MUX21X1 U172(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[3]) ,.Q(int_map_req_v[172]));
	MUX21X1 U173(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[3]) ,.Q(int_map_req_v[173]));
	MUX21X1 U174(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[3]) ,.Q(int_map_req_v[174]));
	MUX21X1 U175(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[3]) ,.Q(int_map_req_v[175]));
	MUX21X1 U176(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[3]) ,.Q(int_map_req_v[176]));
	MUX21X1 U177(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[3]) ,.Q(int_map_req_v[177]));
	MUX21X1 U178(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[3]) ,.Q(int_map_req_v[178]));
	MUX21X1 U179(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[3]) ,.Q(int_map_req_v[179]));
	MUX21X1 U180(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[3]) ,.Q(int_map_req_v[180]));
	MUX21X1 U181(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[3]) ,.Q(int_map_req_v[181]));
	MUX21X1 U182(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[3]) ,.Q(int_map_req_v[182]));
	MUX21X1 U183(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[3]) ,.Q(int_map_req_v[183]));
	MUX21X1 U184(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[3]) ,.Q(int_map_req_v[184]));
	MUX21X1 U185(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[23]) ,.Q(int_map_req_v[185]));
	MUX21X1 U186(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[23]) ,.Q(int_map_req_v[186]));
	MUX21X1 U187(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[23]) ,.Q(int_map_req_v[187]));
	MUX21X1 U188(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[23]) ,.Q(int_map_req_v[188]));
	MUX21X1 U189(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[23]) ,.Q(int_map_req_v[189]));
	MUX21X1 U190(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[23]) ,.Q(int_map_req_v[190]));
	MUX21X1 U191(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[23]) ,.Q(int_map_req_v[191]));
	MUX21X1 U192(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[23]) ,.Q(int_map_req_v[192]));
	MUX21X1 U193(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[23]) ,.Q(int_map_req_v[193]));
	MUX21X1 U194(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[23]) ,.Q(int_map_req_v[194]));
	MUX21X1 U195(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[23]) ,.Q(int_map_req_v[195]));
	MUX21X1 U196(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[23]) ,.Q(int_map_req_v[196]));
	MUX21X1 U197(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[23]) ,.Q(int_map_req_v[197]));
	MUX21X1 U198(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[23]) ,.Q(int_map_req_v[198]));
	MUX21X1 U199(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[23]) ,.Q(int_map_req_v[199]));
	MUX21X1 U200(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[23]) ,.Q(int_map_req_v[200]));
	MUX21X1 U201(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[23]) ,.Q(int_map_req_v[201]));
	MUX21X1 U202(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[23]) ,.Q(int_map_req_v[202]));
	MUX21X1 U203(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[23]) ,.Q(int_map_req_v[203]));
	MUX21X1 U204(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[23]) ,.Q(int_map_req_v[204]));
	MUX21X1 U205(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[23]) ,.Q(int_map_req_v[205]));
	MUX21X1 U206(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[23]) ,.Q(int_map_req_v[206]));
	MUX21X1 U207(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[23]) ,.Q(int_map_req_v[207]));
	MUX21X1 U208(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[23]) ,.Q(int_map_req_v[208]));
	MUX21X1 U209(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[23]) ,.Q(int_map_req_v[209]));
	MUX21X1 U210(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[23]) ,.Q(int_map_req_v[210]));
	MUX21X1 U211(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[23]) ,.Q(int_map_req_v[211]));
	MUX21X1 U212(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[23]) ,.Q(int_map_req_v[212]));
	MUX21X1 U213(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[23]) ,.Q(int_map_req_v[213]));
	MUX21X1 U214(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[23]) ,.Q(int_map_req_v[214]));
	MUX21X1 U215(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[23]) ,.Q(int_map_req_v[215]));
	MUX21X1 U216(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[23]) ,.Q(int_map_req_v[216]));
	MUX21X1 U217(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[23]) ,.Q(int_map_req_v[217]));
	MUX21X1 U218(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[23]) ,.Q(int_map_req_v[218]));
	MUX21X1 U219(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[23]) ,.Q(int_map_req_v[219]));
	MUX21X1 U220(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[23]) ,.Q(int_map_req_v[220]));
	MUX21X1 U221(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[23]) ,.Q(int_map_req_v[221]));
	MUX21X1 U222(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[18]) ,.Q(int_map_req_v[222]));
	MUX21X1 U223(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[18]) ,.Q(int_map_req_v[223]));
	MUX21X1 U224(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[18]) ,.Q(int_map_req_v[224]));
	MUX21X1 U225(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[18]) ,.Q(int_map_req_v[225]));
	MUX21X1 U226(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[18]) ,.Q(int_map_req_v[226]));
	MUX21X1 U227(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[18]) ,.Q(int_map_req_v[227]));
	MUX21X1 U228(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[18]) ,.Q(int_map_req_v[228]));
	MUX21X1 U229(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[18]) ,.Q(int_map_req_v[229]));
	MUX21X1 U230(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[18]) ,.Q(int_map_req_v[230]));
	MUX21X1 U231(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[18]) ,.Q(int_map_req_v[231]));
	MUX21X1 U232(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[18]) ,.Q(int_map_req_v[232]));
	MUX21X1 U233(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[18]) ,.Q(int_map_req_v[233]));
	MUX21X1 U234(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[18]) ,.Q(int_map_req_v[234]));
	MUX21X1 U235(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[18]) ,.Q(int_map_req_v[235]));
	MUX21X1 U236(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[18]) ,.Q(int_map_req_v[236]));
	MUX21X1 U237(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[18]) ,.Q(int_map_req_v[237]));
	MUX21X1 U238(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[18]) ,.Q(int_map_req_v[238]));
	MUX21X1 U239(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[18]) ,.Q(int_map_req_v[239]));
	MUX21X1 U240(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[18]) ,.Q(int_map_req_v[240]));
	MUX21X1 U241(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[18]) ,.Q(int_map_req_v[241]));
	MUX21X1 U242(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[18]) ,.Q(int_map_req_v[242]));
	MUX21X1 U243(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[18]) ,.Q(int_map_req_v[243]));
	MUX21X1 U244(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[18]) ,.Q(int_map_req_v[244]));
	MUX21X1 U245(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[18]) ,.Q(int_map_req_v[245]));
	MUX21X1 U246(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[18]) ,.Q(int_map_req_v[246]));
	MUX21X1 U247(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[18]) ,.Q(int_map_req_v[247]));
	MUX21X1 U248(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[18]) ,.Q(int_map_req_v[248]));
	MUX21X1 U249(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[18]) ,.Q(int_map_req_v[249]));
	MUX21X1 U250(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[18]) ,.Q(int_map_req_v[250]));
	MUX21X1 U251(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[18]) ,.Q(int_map_req_v[251]));
	MUX21X1 U252(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[18]) ,.Q(int_map_req_v[252]));
	MUX21X1 U253(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[18]) ,.Q(int_map_req_v[253]));
	MUX21X1 U254(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[18]) ,.Q(int_map_req_v[254]));
	MUX21X1 U255(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[18]) ,.Q(int_map_req_v[255]));
	MUX21X1 U256(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[18]) ,.Q(int_map_req_v[256]));
	MUX21X1 U257(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[18]) ,.Q(int_map_req_v[257]));
	MUX21X1 U258(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[18]) ,.Q(int_map_req_v[258]));
	MUX21X1 U259(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[13]) ,.Q(int_map_req_v[259]));
	MUX21X1 U260(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[13]) ,.Q(int_map_req_v[260]));
	MUX21X1 U261(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[13]) ,.Q(int_map_req_v[261]));
	MUX21X1 U262(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[13]) ,.Q(int_map_req_v[262]));
	MUX21X1 U263(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[13]) ,.Q(int_map_req_v[263]));
	MUX21X1 U264(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[13]) ,.Q(int_map_req_v[264]));
	MUX21X1 U265(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[13]) ,.Q(int_map_req_v[265]));
	MUX21X1 U266(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[13]) ,.Q(int_map_req_v[266]));
	MUX21X1 U267(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[13]) ,.Q(int_map_req_v[267]));
	MUX21X1 U268(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[13]) ,.Q(int_map_req_v[268]));
	MUX21X1 U269(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[13]) ,.Q(int_map_req_v[269]));
	MUX21X1 U270(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[13]) ,.Q(int_map_req_v[270]));
	MUX21X1 U271(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[13]) ,.Q(int_map_req_v[271]));
	MUX21X1 U272(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[13]) ,.Q(int_map_req_v[272]));
	MUX21X1 U273(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[13]) ,.Q(int_map_req_v[273]));
	MUX21X1 U274(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[13]) ,.Q(int_map_req_v[274]));
	MUX21X1 U275(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[13]) ,.Q(int_map_req_v[275]));
	MUX21X1 U276(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[13]) ,.Q(int_map_req_v[276]));
	MUX21X1 U277(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[13]) ,.Q(int_map_req_v[277]));
	MUX21X1 U278(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[13]) ,.Q(int_map_req_v[278]));
	MUX21X1 U279(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[13]) ,.Q(int_map_req_v[279]));
	MUX21X1 U280(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[13]) ,.Q(int_map_req_v[280]));
	MUX21X1 U281(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[13]) ,.Q(int_map_req_v[281]));
	MUX21X1 U282(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[13]) ,.Q(int_map_req_v[282]));
	MUX21X1 U283(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[13]) ,.Q(int_map_req_v[283]));
	MUX21X1 U284(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[13]) ,.Q(int_map_req_v[284]));
	MUX21X1 U285(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[13]) ,.Q(int_map_req_v[285]));
	MUX21X1 U286(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[13]) ,.Q(int_map_req_v[286]));
	MUX21X1 U287(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[13]) ,.Q(int_map_req_v[287]));
	MUX21X1 U288(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[13]) ,.Q(int_map_req_v[288]));
	MUX21X1 U289(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[13]) ,.Q(int_map_req_v[289]));
	MUX21X1 U290(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[13]) ,.Q(int_map_req_v[290]));
	MUX21X1 U291(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[13]) ,.Q(int_map_req_v[291]));
	MUX21X1 U292(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[13]) ,.Q(int_map_req_v[292]));
	MUX21X1 U293(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[13]) ,.Q(int_map_req_v[293]));
	MUX21X1 U294(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[13]) ,.Q(int_map_req_v[294]));
	MUX21X1 U295(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[13]) ,.Q(int_map_req_v[295]));
	MUX21X1 U09(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[7]), .S(int_route_v[13]) ,.Q(int_resp_v[2]));
	MUX21X1 U10(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[8]), .S(int_route_v[13]) ,.Q(int_resp_v[3]));
	MUX21X1 U11(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[6]), .S(int_route_v[18]) ,.Q(int_resp_v[3]));
	MUX21X1 U12(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[7]), .S(int_route_v[18]) ,.Q(int_resp_v[4]));
	MUX21X1 U13(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[4]));
	MUX21X1 U14(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[2]), .S(int_route_v[6]) ,.Q(int_resp_v[5]));
	MUX21X1 U15(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[0]), .S(int_route_v[4]) ,.Q(int_resp_v[0]));
	MUX21X1 U16(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));


	MUX21X1 U296(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[7]) ,.Q(int_map_req_v[296]));
	MUX21X1 U297(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[7]) ,.Q(int_map_req_v[297]));
	MUX21X1 U298(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[7]) ,.Q(int_map_req_v[298]));
	MUX21X1 U299(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[7]) ,.Q(int_map_req_v[299]));
	MUX21X1 U300(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[7]) ,.Q(int_map_req_v[300]));
	MUX21X1 U301(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[7]) ,.Q(int_map_req_v[301]));
	MUX21X1 U302(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[7]) ,.Q(int_map_req_v[302]));
	MUX21X1 U303(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[7]) ,.Q(int_map_req_v[303]));
	MUX21X1 U304(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[7]) ,.Q(int_map_req_v[304]));
	MUX21X1 U305(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[7]) ,.Q(int_map_req_v[305]));
	MUX21X1 U306(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[7]) ,.Q(int_map_req_v[306]));
	MUX21X1 U307(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[7]) ,.Q(int_map_req_v[307]));
	MUX21X1 U308(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[7]) ,.Q(int_map_req_v[308]));
	MUX21X1 U309(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[7]) ,.Q(int_map_req_v[309]));
	MUX21X1 U310(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[7]) ,.Q(int_map_req_v[310]));
	MUX21X1 U311(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[7]) ,.Q(int_map_req_v[311]));
	MUX21X1 U312(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[7]) ,.Q(int_map_req_v[312]));
	MUX21X1 U313(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[7]) ,.Q(int_map_req_v[313]));
	MUX21X1 U314(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[7]) ,.Q(int_map_req_v[314]));
	MUX21X1 U315(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[7]) ,.Q(int_map_req_v[315]));
	MUX21X1 U316(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[7]) ,.Q(int_map_req_v[316]));
	MUX21X1 U317(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[7]) ,.Q(int_map_req_v[317]));
	MUX21X1 U318(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[7]) ,.Q(int_map_req_v[318]));
	MUX21X1 U319(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[7]) ,.Q(int_map_req_v[319]));
	MUX21X1 U320(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[7]) ,.Q(int_map_req_v[320]));
	MUX21X1 U321(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[7]) ,.Q(int_map_req_v[321]));
	MUX21X1 U322(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[7]) ,.Q(int_map_req_v[322]));
	MUX21X1 U323(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[7]) ,.Q(int_map_req_v[323]));
	MUX21X1 U324(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[7]) ,.Q(int_map_req_v[324]));
	MUX21X1 U325(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[7]) ,.Q(int_map_req_v[325]));
	MUX21X1 U326(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[7]) ,.Q(int_map_req_v[326]));
	MUX21X1 U327(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[7]) ,.Q(int_map_req_v[327]));
	MUX21X1 U328(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[7]) ,.Q(int_map_req_v[328]));
	MUX21X1 U329(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[7]) ,.Q(int_map_req_v[329]));
	MUX21X1 U330(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[7]) ,.Q(int_map_req_v[330]));
	MUX21X1 U331(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[7]) ,.Q(int_map_req_v[331]));
	MUX21X1 U332(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[7]) ,.Q(int_map_req_v[332]));
	MUX21X1 U333(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[2]) ,.Q(int_map_req_v[333]));
	MUX21X1 U334(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[2]) ,.Q(int_map_req_v[334]));
	MUX21X1 U335(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[2]) ,.Q(int_map_req_v[335]));
	MUX21X1 U336(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[2]) ,.Q(int_map_req_v[336]));
	MUX21X1 U337(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[2]) ,.Q(int_map_req_v[337]));
	MUX21X1 U338(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[2]) ,.Q(int_map_req_v[338]));
	MUX21X1 U339(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[2]) ,.Q(int_map_req_v[339]));
	MUX21X1 U340(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[2]) ,.Q(int_map_req_v[340]));
	MUX21X1 U341(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[2]) ,.Q(int_map_req_v[341]));
	MUX21X1 U342(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[2]) ,.Q(int_map_req_v[342]));
	MUX21X1 U343(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[2]) ,.Q(int_map_req_v[343]));
	MUX21X1 U344(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[2]) ,.Q(int_map_req_v[344]));
	MUX21X1 U345(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[2]) ,.Q(int_map_req_v[345]));
	MUX21X1 U346(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[2]) ,.Q(int_map_req_v[346]));
	MUX21X1 U347(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[2]) ,.Q(int_map_req_v[347]));
	MUX21X1 U348(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[2]) ,.Q(int_map_req_v[348]));
	MUX21X1 U349(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[2]) ,.Q(int_map_req_v[349]));
	MUX21X1 U350(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[2]) ,.Q(int_map_req_v[350]));
	MUX21X1 U351(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[2]) ,.Q(int_map_req_v[351]));
	MUX21X1 U352(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[2]) ,.Q(int_map_req_v[352]));
	MUX21X1 U353(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[2]) ,.Q(int_map_req_v[353]));
	MUX21X1 U354(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[2]) ,.Q(int_map_req_v[354]));
	MUX21X1 U355(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[2]) ,.Q(int_map_req_v[355]));
	MUX21X1 U356(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[2]) ,.Q(int_map_req_v[356]));
	MUX21X1 U357(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[2]) ,.Q(int_map_req_v[357]));
	MUX21X1 U358(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[2]) ,.Q(int_map_req_v[358]));
	MUX21X1 U359(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[2]) ,.Q(int_map_req_v[359]));
	MUX21X1 U360(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[2]) ,.Q(int_map_req_v[360]));
	MUX21X1 U361(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[2]) ,.Q(int_map_req_v[361]));
	MUX21X1 U362(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[2]) ,.Q(int_map_req_v[362]));
	MUX21X1 U363(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[2]) ,.Q(int_map_req_v[363]));
	MUX21X1 U364(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[2]) ,.Q(int_map_req_v[364]));
	MUX21X1 U365(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[2]) ,.Q(int_map_req_v[365]));
	MUX21X1 U366(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[2]) ,.Q(int_map_req_v[366]));
	MUX21X1 U367(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[2]) ,.Q(int_map_req_v[367]));
	MUX21X1 U368(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[2]) ,.Q(int_map_req_v[368]));
	MUX21X1 U369(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[2]) ,.Q(int_map_req_v[369]));
	MUX21X1 U370(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[22]) ,.Q(int_map_req_v[370]));
	MUX21X1 U371(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[22]) ,.Q(int_map_req_v[371]));
	MUX21X1 U372(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[22]) ,.Q(int_map_req_v[372]));
	MUX21X1 U373(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[22]) ,.Q(int_map_req_v[373]));
	MUX21X1 U374(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[22]) ,.Q(int_map_req_v[374]));
	MUX21X1 U375(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[22]) ,.Q(int_map_req_v[375]));
	MUX21X1 U376(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[22]) ,.Q(int_map_req_v[376]));
	MUX21X1 U377(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[22]) ,.Q(int_map_req_v[377]));
	MUX21X1 U378(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[22]) ,.Q(int_map_req_v[378]));
	MUX21X1 U379(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[22]) ,.Q(int_map_req_v[379]));
	MUX21X1 U380(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[22]) ,.Q(int_map_req_v[380]));
	MUX21X1 U381(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[22]) ,.Q(int_map_req_v[381]));
	MUX21X1 U382(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[22]) ,.Q(int_map_req_v[382]));
	MUX21X1 U383(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[22]) ,.Q(int_map_req_v[383]));
	MUX21X1 U384(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[22]) ,.Q(int_map_req_v[384]));
	MUX21X1 U385(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[22]) ,.Q(int_map_req_v[385]));
	MUX21X1 U386(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[22]) ,.Q(int_map_req_v[386]));
	MUX21X1 U387(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[22]) ,.Q(int_map_req_v[387]));
	MUX21X1 U388(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[22]) ,.Q(int_map_req_v[388]));
	MUX21X1 U389(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[22]) ,.Q(int_map_req_v[389]));
	MUX21X1 U390(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[22]) ,.Q(int_map_req_v[390]));
	MUX21X1 U391(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[22]) ,.Q(int_map_req_v[391]));
	MUX21X1 U392(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[22]) ,.Q(int_map_req_v[392]));
	MUX21X1 U393(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[22]) ,.Q(int_map_req_v[393]));
	MUX21X1 U394(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[22]) ,.Q(int_map_req_v[394]));
	MUX21X1 U395(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[22]) ,.Q(int_map_req_v[395]));
	MUX21X1 U396(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[22]) ,.Q(int_map_req_v[396]));
	MUX21X1 U397(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[22]) ,.Q(int_map_req_v[397]));
	MUX21X1 U398(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[22]) ,.Q(int_map_req_v[398]));
	MUX21X1 U399(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[22]) ,.Q(int_map_req_v[399]));
	MUX21X1 U400(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[22]) ,.Q(int_map_req_v[400]));
	MUX21X1 U401(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[22]) ,.Q(int_map_req_v[401]));
	MUX21X1 U402(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[22]) ,.Q(int_map_req_v[402]));
	MUX21X1 U403(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[22]) ,.Q(int_map_req_v[403]));
	MUX21X1 U404(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[22]) ,.Q(int_map_req_v[404]));
	MUX21X1 U405(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[22]) ,.Q(int_map_req_v[405]));
	MUX21X1 U406(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[22]) ,.Q(int_map_req_v[406]));
	MUX21X1 U407(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[17]) ,.Q(int_map_req_v[407]));
	MUX21X1 U408(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[17]) ,.Q(int_map_req_v[408]));
	MUX21X1 U409(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[17]) ,.Q(int_map_req_v[409]));
	MUX21X1 U410(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[17]) ,.Q(int_map_req_v[410]));
	MUX21X1 U411(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[17]) ,.Q(int_map_req_v[411]));
	MUX21X1 U412(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[17]) ,.Q(int_map_req_v[412]));
	MUX21X1 U413(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[17]) ,.Q(int_map_req_v[413]));
	MUX21X1 U414(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[17]) ,.Q(int_map_req_v[414]));
	MUX21X1 U415(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[17]) ,.Q(int_map_req_v[415]));
	MUX21X1 U416(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[17]) ,.Q(int_map_req_v[416]));
	MUX21X1 U417(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[17]) ,.Q(int_map_req_v[417]));
	MUX21X1 U418(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[17]) ,.Q(int_map_req_v[418]));
	MUX21X1 U419(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[17]) ,.Q(int_map_req_v[419]));
	MUX21X1 U420(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[17]) ,.Q(int_map_req_v[420]));
	MUX21X1 U421(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[17]) ,.Q(int_map_req_v[421]));
	MUX21X1 U422(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[17]) ,.Q(int_map_req_v[422]));
	MUX21X1 U423(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[17]) ,.Q(int_map_req_v[423]));
	MUX21X1 U424(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[17]) ,.Q(int_map_req_v[424]));
	MUX21X1 U425(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[17]) ,.Q(int_map_req_v[425]));
	MUX21X1 U426(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[17]) ,.Q(int_map_req_v[426]));
	MUX21X1 U427(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[17]) ,.Q(int_map_req_v[427]));
	MUX21X1 U428(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[17]) ,.Q(int_map_req_v[428]));
	MUX21X1 U429(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[17]) ,.Q(int_map_req_v[429]));
	MUX21X1 U430(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[17]) ,.Q(int_map_req_v[430]));
	MUX21X1 U431(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[17]) ,.Q(int_map_req_v[431]));
	MUX21X1 U432(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[17]) ,.Q(int_map_req_v[432]));
	MUX21X1 U433(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[17]) ,.Q(int_map_req_v[433]));
	MUX21X1 U434(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[17]) ,.Q(int_map_req_v[434]));
	MUX21X1 U435(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[17]) ,.Q(int_map_req_v[435]));
	MUX21X1 U436(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[17]) ,.Q(int_map_req_v[436]));
	MUX21X1 U437(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[17]) ,.Q(int_map_req_v[437]));
	MUX21X1 U438(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[17]) ,.Q(int_map_req_v[438]));
	MUX21X1 U439(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[17]) ,.Q(int_map_req_v[439]));
	MUX21X1 U440(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[17]) ,.Q(int_map_req_v[440]));
	MUX21X1 U441(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[17]) ,.Q(int_map_req_v[441]));
	MUX21X1 U442(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[17]) ,.Q(int_map_req_v[442]));
	MUX21X1 U443(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[17]) ,.Q(int_map_req_v[443]));
	MUX21X1 U17(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[11]), .S(int_route_v[17]) ,.Q(int_resp_v[3]));
	MUX21X1 U18(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[12]), .S(int_route_v[17]) ,.Q(int_resp_v[4]));
	MUX21X1 U19(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[10]), .S(int_route_v[22]) ,.Q(int_resp_v[4]));
	MUX21X1 U20(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[11]), .S(int_route_v[22]) ,.Q(int_resp_v[5]));
	MUX21X1 U21(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[9]), .S(int_route_v[2]) ,.Q(int_resp_v[0]));
	MUX21X1 U22(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[10]), .S(int_route_v[2]) ,.Q(int_resp_v[1]));
	MUX21X1 U23(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[8]), .S(int_route_v[7]) ,.Q(int_resp_v[1]));
	MUX21X1 U24(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[9]), .S(int_route_v[7]) ,.Q(int_resp_v[2]));

	MUX21X1 U444(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[11]) ,.Q(int_map_req_v[444]));
	MUX21X1 U445(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[11]) ,.Q(int_map_req_v[445]));
	MUX21X1 U446(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[11]) ,.Q(int_map_req_v[446]));
	MUX21X1 U447(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[11]) ,.Q(int_map_req_v[447]));
	MUX21X1 U448(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[11]) ,.Q(int_map_req_v[448]));
	MUX21X1 U449(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[11]) ,.Q(int_map_req_v[449]));
	MUX21X1 U450(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[11]) ,.Q(int_map_req_v[450]));
	MUX21X1 U451(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[11]) ,.Q(int_map_req_v[451]));
	MUX21X1 U452(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[11]) ,.Q(int_map_req_v[452]));
	MUX21X1 U453(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[11]) ,.Q(int_map_req_v[453]));
	MUX21X1 U454(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[11]) ,.Q(int_map_req_v[454]));
	MUX21X1 U455(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[11]) ,.Q(int_map_req_v[455]));
	MUX21X1 U456(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[11]) ,.Q(int_map_req_v[456]));
	MUX21X1 U457(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[11]) ,.Q(int_map_req_v[457]));
	MUX21X1 U458(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[11]) ,.Q(int_map_req_v[458]));
	MUX21X1 U459(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[11]) ,.Q(int_map_req_v[459]));
	MUX21X1 U460(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[11]) ,.Q(int_map_req_v[460]));
	MUX21X1 U461(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[11]) ,.Q(int_map_req_v[461]));
	MUX21X1 U462(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[11]) ,.Q(int_map_req_v[462]));
	MUX21X1 U463(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[11]) ,.Q(int_map_req_v[463]));
	MUX21X1 U464(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[11]) ,.Q(int_map_req_v[464]));
	MUX21X1 U465(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[11]) ,.Q(int_map_req_v[465]));
	MUX21X1 U466(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[11]) ,.Q(int_map_req_v[466]));
	MUX21X1 U467(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[11]) ,.Q(int_map_req_v[467]));
	MUX21X1 U468(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[11]) ,.Q(int_map_req_v[468]));
	MUX21X1 U469(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[11]) ,.Q(int_map_req_v[469]));
	MUX21X1 U470(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[11]) ,.Q(int_map_req_v[470]));
	MUX21X1 U471(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[11]) ,.Q(int_map_req_v[471]));
	MUX21X1 U472(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[11]) ,.Q(int_map_req_v[472]));
	MUX21X1 U473(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[11]) ,.Q(int_map_req_v[473]));
	MUX21X1 U474(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[11]) ,.Q(int_map_req_v[474]));
	MUX21X1 U475(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[11]) ,.Q(int_map_req_v[475]));
	MUX21X1 U476(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[11]) ,.Q(int_map_req_v[476]));
	MUX21X1 U477(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[11]) ,.Q(int_map_req_v[477]));
	MUX21X1 U478(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[11]) ,.Q(int_map_req_v[478]));
	MUX21X1 U479(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[11]) ,.Q(int_map_req_v[479]));
	MUX21X1 U480(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[11]) ,.Q(int_map_req_v[480]));
	MUX21X1 U481(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[6]) ,.Q(int_map_req_v[481]));
	MUX21X1 U482(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[6]) ,.Q(int_map_req_v[482]));
	MUX21X1 U483(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[6]) ,.Q(int_map_req_v[483]));
	MUX21X1 U484(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[6]) ,.Q(int_map_req_v[484]));
	MUX21X1 U485(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[6]) ,.Q(int_map_req_v[485]));
	MUX21X1 U486(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[6]) ,.Q(int_map_req_v[486]));
	MUX21X1 U487(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[6]) ,.Q(int_map_req_v[487]));
	MUX21X1 U488(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[6]) ,.Q(int_map_req_v[488]));
	MUX21X1 U489(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[6]) ,.Q(int_map_req_v[489]));
	MUX21X1 U490(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[6]) ,.Q(int_map_req_v[490]));
	MUX21X1 U491(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[6]) ,.Q(int_map_req_v[491]));
	MUX21X1 U492(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[6]) ,.Q(int_map_req_v[492]));
	MUX21X1 U493(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[6]) ,.Q(int_map_req_v[493]));
	MUX21X1 U494(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[6]) ,.Q(int_map_req_v[494]));
	MUX21X1 U495(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[6]) ,.Q(int_map_req_v[495]));
	MUX21X1 U496(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[6]) ,.Q(int_map_req_v[496]));
	MUX21X1 U497(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[6]) ,.Q(int_map_req_v[497]));
	MUX21X1 U498(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[6]) ,.Q(int_map_req_v[498]));
	MUX21X1 U499(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[6]) ,.Q(int_map_req_v[499]));
	MUX21X1 U500(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[6]) ,.Q(int_map_req_v[500]));
	MUX21X1 U501(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[6]) ,.Q(int_map_req_v[501]));
	MUX21X1 U502(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[6]) ,.Q(int_map_req_v[502]));
	MUX21X1 U503(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[6]) ,.Q(int_map_req_v[503]));
	MUX21X1 U504(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[6]) ,.Q(int_map_req_v[504]));
	MUX21X1 U505(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[6]) ,.Q(int_map_req_v[505]));
	MUX21X1 U506(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[6]) ,.Q(int_map_req_v[506]));
	MUX21X1 U507(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[6]) ,.Q(int_map_req_v[507]));
	MUX21X1 U508(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[6]) ,.Q(int_map_req_v[508]));
	MUX21X1 U509(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[6]) ,.Q(int_map_req_v[509]));
	MUX21X1 U510(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[6]) ,.Q(int_map_req_v[510]));
	MUX21X1 U511(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[6]) ,.Q(int_map_req_v[511]));
	MUX21X1 U512(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[6]) ,.Q(int_map_req_v[512]));
	MUX21X1 U513(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[6]) ,.Q(int_map_req_v[513]));
	MUX21X1 U514(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[6]) ,.Q(int_map_req_v[514]));
	MUX21X1 U515(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[6]) ,.Q(int_map_req_v[515]));
	MUX21X1 U516(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[6]) ,.Q(int_map_req_v[516]));
	MUX21X1 U517(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[6]) ,.Q(int_map_req_v[517]));
	MUX21X1 U518(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[1]) ,.Q(int_map_req_v[518]));
	MUX21X1 U519(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[1]) ,.Q(int_map_req_v[519]));
	MUX21X1 U520(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[1]) ,.Q(int_map_req_v[520]));
	MUX21X1 U521(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[1]) ,.Q(int_map_req_v[521]));
	MUX21X1 U522(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[1]) ,.Q(int_map_req_v[522]));
	MUX21X1 U523(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[1]) ,.Q(int_map_req_v[523]));
	MUX21X1 U524(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[1]) ,.Q(int_map_req_v[524]));
	MUX21X1 U525(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[1]) ,.Q(int_map_req_v[525]));
	MUX21X1 U526(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[1]) ,.Q(int_map_req_v[526]));
	MUX21X1 U527(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[1]) ,.Q(int_map_req_v[527]));
	MUX21X1 U528(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[1]) ,.Q(int_map_req_v[528]));
	MUX21X1 U529(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[1]) ,.Q(int_map_req_v[529]));
	MUX21X1 U530(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[1]) ,.Q(int_map_req_v[530]));
	MUX21X1 U531(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[1]) ,.Q(int_map_req_v[531]));
	MUX21X1 U532(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[1]) ,.Q(int_map_req_v[532]));
	MUX21X1 U533(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[1]) ,.Q(int_map_req_v[533]));
	MUX21X1 U534(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[1]) ,.Q(int_map_req_v[534]));
	MUX21X1 U535(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[1]) ,.Q(int_map_req_v[535]));
	MUX21X1 U536(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[1]) ,.Q(int_map_req_v[536]));
	MUX21X1 U537(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[1]) ,.Q(int_map_req_v[537]));
	MUX21X1 U538(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[1]) ,.Q(int_map_req_v[538]));
	MUX21X1 U539(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[1]) ,.Q(int_map_req_v[539]));
	MUX21X1 U540(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[1]) ,.Q(int_map_req_v[540]));
	MUX21X1 U541(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[1]) ,.Q(int_map_req_v[541]));
	MUX21X1 U542(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[1]) ,.Q(int_map_req_v[542]));
	MUX21X1 U543(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[1]) ,.Q(int_map_req_v[543]));
	MUX21X1 U544(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[1]) ,.Q(int_map_req_v[544]));
	MUX21X1 U545(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[1]) ,.Q(int_map_req_v[545]));
	MUX21X1 U546(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[1]) ,.Q(int_map_req_v[546]));
	MUX21X1 U547(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[1]) ,.Q(int_map_req_v[547]));
	MUX21X1 U548(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[1]) ,.Q(int_map_req_v[548]));
	MUX21X1 U549(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[1]) ,.Q(int_map_req_v[549]));
	MUX21X1 U550(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[1]) ,.Q(int_map_req_v[550]));
	MUX21X1 U551(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[1]) ,.Q(int_map_req_v[551]));
	MUX21X1 U552(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[1]) ,.Q(int_map_req_v[552]));
	MUX21X1 U553(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[1]) ,.Q(int_map_req_v[553]));
	MUX21X1 U554(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[1]) ,.Q(int_map_req_v[554]));
	MUX21X1 U555(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[21]) ,.Q(int_map_req_v[555]));
	MUX21X1 U556(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[21]) ,.Q(int_map_req_v[556]));
	MUX21X1 U557(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[21]) ,.Q(int_map_req_v[557]));
	MUX21X1 U558(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[21]) ,.Q(int_map_req_v[558]));
	MUX21X1 U559(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[21]) ,.Q(int_map_req_v[559]));
	MUX21X1 U560(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[21]) ,.Q(int_map_req_v[560]));
	MUX21X1 U561(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[21]) ,.Q(int_map_req_v[561]));
	MUX21X1 U562(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[21]) ,.Q(int_map_req_v[562]));
	MUX21X1 U563(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[21]) ,.Q(int_map_req_v[563]));
	MUX21X1 U564(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[21]) ,.Q(int_map_req_v[564]));
	MUX21X1 U565(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[21]) ,.Q(int_map_req_v[565]));
	MUX21X1 U566(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[21]) ,.Q(int_map_req_v[566]));
	MUX21X1 U567(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[21]) ,.Q(int_map_req_v[567]));
	MUX21X1 U568(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[21]) ,.Q(int_map_req_v[568]));
	MUX21X1 U569(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[21]) ,.Q(int_map_req_v[569]));
	MUX21X1 U570(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[21]) ,.Q(int_map_req_v[570]));
	MUX21X1 U571(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[21]) ,.Q(int_map_req_v[571]));
	MUX21X1 U572(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[21]) ,.Q(int_map_req_v[572]));
	MUX21X1 U573(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[21]) ,.Q(int_map_req_v[573]));
	MUX21X1 U574(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[21]) ,.Q(int_map_req_v[574]));
	MUX21X1 U575(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[21]) ,.Q(int_map_req_v[575]));
	MUX21X1 U576(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[21]) ,.Q(int_map_req_v[576]));
	MUX21X1 U577(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[21]) ,.Q(int_map_req_v[577]));
	MUX21X1 U578(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[21]) ,.Q(int_map_req_v[578]));
	MUX21X1 U579(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[21]) ,.Q(int_map_req_v[579]));
	MUX21X1 U580(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[21]) ,.Q(int_map_req_v[580]));
	MUX21X1 U581(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[21]) ,.Q(int_map_req_v[581]));
	MUX21X1 U582(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[21]) ,.Q(int_map_req_v[582]));
	MUX21X1 U583(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[21]) ,.Q(int_map_req_v[583]));
	MUX21X1 U584(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[21]) ,.Q(int_map_req_v[584]));
	MUX21X1 U585(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[21]) ,.Q(int_map_req_v[585]));
	MUX21X1 U586(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[21]) ,.Q(int_map_req_v[586]));
	MUX21X1 U587(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[21]) ,.Q(int_map_req_v[587]));
	MUX21X1 U588(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[21]) ,.Q(int_map_req_v[588]));
	MUX21X1 U589(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[21]) ,.Q(int_map_req_v[589]));
	MUX21X1 U590(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[21]) ,.Q(int_map_req_v[590]));
	MUX21X1 U591(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[21]) ,.Q(int_map_req_v[591]));
	MUX21X1 U25(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[15]), .S(int_route_v[21]) ,.Q(int_resp_v[4]));
	MUX21X1 U26(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[16]), .S(int_route_v[21]) ,.Q(int_resp_v[5]));
	MUX21X1 U27(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[14]), .S(int_route_v[1]) ,.Q(int_resp_v[0]));
	MUX21X1 U28(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[15]), .S(int_route_v[1]) ,.Q(int_resp_v[1]));
	MUX21X1 U29(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[13]), .S(int_route_v[6]) ,.Q(int_resp_v[1]));
	MUX21X1 U30(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[14]), .S(int_route_v[6]) ,.Q(int_resp_v[2]));
	MUX21X1 U31(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[12]), .S(int_route_v[11]) ,.Q(int_resp_v[2]));
	MUX21X1 U32(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[13]), .S(int_route_v[11]) ,.Q(int_resp_v[3]));



	MUX21X1 U592(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[15]) ,.Q(int_map_req_v[592]));
	MUX21X1 U593(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[15]) ,.Q(int_map_req_v[593]));
	MUX21X1 U594(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[15]) ,.Q(int_map_req_v[594]));
	MUX21X1 U595(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[15]) ,.Q(int_map_req_v[595]));
	MUX21X1 U596(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[15]) ,.Q(int_map_req_v[596]));
	MUX21X1 U597(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[15]) ,.Q(int_map_req_v[597]));
	MUX21X1 U598(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[15]) ,.Q(int_map_req_v[598]));
	MUX21X1 U599(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[15]) ,.Q(int_map_req_v[599]));
	MUX21X1 U600(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[15]) ,.Q(int_map_req_v[600]));
	MUX21X1 U601(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[15]) ,.Q(int_map_req_v[601]));
	MUX21X1 U602(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[15]) ,.Q(int_map_req_v[602]));
	MUX21X1 U603(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[15]) ,.Q(int_map_req_v[603]));
	MUX21X1 U604(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[15]) ,.Q(int_map_req_v[604]));
	MUX21X1 U605(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[15]) ,.Q(int_map_req_v[605]));
	MUX21X1 U606(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[15]) ,.Q(int_map_req_v[606]));
	MUX21X1 U607(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[15]) ,.Q(int_map_req_v[607]));
	MUX21X1 U608(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[15]) ,.Q(int_map_req_v[608]));
	MUX21X1 U609(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[15]) ,.Q(int_map_req_v[609]));
	MUX21X1 U610(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[15]) ,.Q(int_map_req_v[610]));
	MUX21X1 U611(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[15]) ,.Q(int_map_req_v[611]));
	MUX21X1 U612(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[15]) ,.Q(int_map_req_v[612]));
	MUX21X1 U613(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[15]) ,.Q(int_map_req_v[613]));
	MUX21X1 U614(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[15]) ,.Q(int_map_req_v[614]));
	MUX21X1 U615(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[15]) ,.Q(int_map_req_v[615]));
	MUX21X1 U616(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[15]) ,.Q(int_map_req_v[616]));
	MUX21X1 U617(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[15]) ,.Q(int_map_req_v[617]));
	MUX21X1 U618(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[15]) ,.Q(int_map_req_v[618]));
	MUX21X1 U619(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[15]) ,.Q(int_map_req_v[619]));
	MUX21X1 U620(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[15]) ,.Q(int_map_req_v[620]));
	MUX21X1 U621(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[15]) ,.Q(int_map_req_v[621]));
	MUX21X1 U622(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[15]) ,.Q(int_map_req_v[622]));
	MUX21X1 U623(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[15]) ,.Q(int_map_req_v[623]));
	MUX21X1 U624(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[15]) ,.Q(int_map_req_v[624]));
	MUX21X1 U625(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[15]) ,.Q(int_map_req_v[625]));
	MUX21X1 U626(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[15]) ,.Q(int_map_req_v[626]));
	MUX21X1 U627(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[15]) ,.Q(int_map_req_v[627]));
	MUX21X1 U628(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[15]) ,.Q(int_map_req_v[628]));
	MUX21X1 U629(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[10]) ,.Q(int_map_req_v[629]));
	MUX21X1 U630(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[10]) ,.Q(int_map_req_v[630]));
	MUX21X1 U631(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[10]) ,.Q(int_map_req_v[631]));
	MUX21X1 U632(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[10]) ,.Q(int_map_req_v[632]));
	MUX21X1 U633(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[10]) ,.Q(int_map_req_v[633]));
	MUX21X1 U634(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[10]) ,.Q(int_map_req_v[634]));
	MUX21X1 U635(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[10]) ,.Q(int_map_req_v[635]));
	MUX21X1 U636(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[10]) ,.Q(int_map_req_v[636]));
	MUX21X1 U637(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[10]) ,.Q(int_map_req_v[637]));
	MUX21X1 U638(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[10]) ,.Q(int_map_req_v[638]));
	MUX21X1 U639(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[10]) ,.Q(int_map_req_v[639]));
	MUX21X1 U640(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[10]) ,.Q(int_map_req_v[640]));
	MUX21X1 U641(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[10]) ,.Q(int_map_req_v[641]));
	MUX21X1 U642(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[10]) ,.Q(int_map_req_v[642]));
	MUX21X1 U643(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[10]) ,.Q(int_map_req_v[643]));
	MUX21X1 U644(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[10]) ,.Q(int_map_req_v[644]));
	MUX21X1 U645(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[10]) ,.Q(int_map_req_v[645]));
	MUX21X1 U646(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[10]) ,.Q(int_map_req_v[646]));
	MUX21X1 U647(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[10]) ,.Q(int_map_req_v[647]));
	MUX21X1 U648(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[10]) ,.Q(int_map_req_v[648]));
	MUX21X1 U649(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[10]) ,.Q(int_map_req_v[649]));
	MUX21X1 U650(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[10]) ,.Q(int_map_req_v[650]));
	MUX21X1 U651(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[10]) ,.Q(int_map_req_v[651]));
	MUX21X1 U652(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[10]) ,.Q(int_map_req_v[652]));
	MUX21X1 U653(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[10]) ,.Q(int_map_req_v[653]));
	MUX21X1 U654(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[10]) ,.Q(int_map_req_v[654]));
	MUX21X1 U655(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[10]) ,.Q(int_map_req_v[655]));
	MUX21X1 U656(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[10]) ,.Q(int_map_req_v[656]));
	MUX21X1 U657(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[10]) ,.Q(int_map_req_v[657]));
	MUX21X1 U658(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[10]) ,.Q(int_map_req_v[658]));
	MUX21X1 U659(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[10]) ,.Q(int_map_req_v[659]));
	MUX21X1 U660(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[10]) ,.Q(int_map_req_v[660]));
	MUX21X1 U661(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[10]) ,.Q(int_map_req_v[661]));
	MUX21X1 U662(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[10]) ,.Q(int_map_req_v[662]));
	MUX21X1 U663(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[10]) ,.Q(int_map_req_v[663]));
	MUX21X1 U664(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[10]) ,.Q(int_map_req_v[664]));
	MUX21X1 U665(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[10]) ,.Q(int_map_req_v[665]));
	MUX21X1 U666(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[5]) ,.Q(int_map_req_v[666]));
	MUX21X1 U667(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[5]) ,.Q(int_map_req_v[667]));
	MUX21X1 U668(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[5]) ,.Q(int_map_req_v[668]));
	MUX21X1 U669(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[5]) ,.Q(int_map_req_v[669]));
	MUX21X1 U670(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[5]) ,.Q(int_map_req_v[670]));
	MUX21X1 U671(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[5]) ,.Q(int_map_req_v[671]));
	MUX21X1 U672(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[5]) ,.Q(int_map_req_v[672]));
	MUX21X1 U673(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[5]) ,.Q(int_map_req_v[673]));
	MUX21X1 U674(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[5]) ,.Q(int_map_req_v[674]));
	MUX21X1 U675(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[5]) ,.Q(int_map_req_v[675]));
	MUX21X1 U676(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[5]) ,.Q(int_map_req_v[676]));
	MUX21X1 U677(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[5]) ,.Q(int_map_req_v[677]));
	MUX21X1 U678(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[5]) ,.Q(int_map_req_v[678]));
	MUX21X1 U679(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[5]) ,.Q(int_map_req_v[679]));
	MUX21X1 U680(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[5]) ,.Q(int_map_req_v[680]));
	MUX21X1 U681(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[5]) ,.Q(int_map_req_v[681]));
	MUX21X1 U682(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[5]) ,.Q(int_map_req_v[682]));
	MUX21X1 U683(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[5]) ,.Q(int_map_req_v[683]));
	MUX21X1 U684(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[5]) ,.Q(int_map_req_v[684]));
	MUX21X1 U685(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[5]) ,.Q(int_map_req_v[685]));
	MUX21X1 U686(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[5]) ,.Q(int_map_req_v[686]));
	MUX21X1 U687(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[5]) ,.Q(int_map_req_v[687]));
	MUX21X1 U688(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[5]) ,.Q(int_map_req_v[688]));
	MUX21X1 U689(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[5]) ,.Q(int_map_req_v[689]));
	MUX21X1 U690(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[5]) ,.Q(int_map_req_v[690]));
	MUX21X1 U691(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[5]) ,.Q(int_map_req_v[691]));
	MUX21X1 U692(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[5]) ,.Q(int_map_req_v[692]));
	MUX21X1 U693(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[5]) ,.Q(int_map_req_v[693]));
	MUX21X1 U694(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[5]) ,.Q(int_map_req_v[694]));
	MUX21X1 U695(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[5]) ,.Q(int_map_req_v[695]));
	MUX21X1 U696(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[5]) ,.Q(int_map_req_v[696]));
	MUX21X1 U697(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[5]) ,.Q(int_map_req_v[697]));
	MUX21X1 U698(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[5]) ,.Q(int_map_req_v[698]));
	MUX21X1 U699(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[5]) ,.Q(int_map_req_v[699]));
	MUX21X1 U700(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[5]) ,.Q(int_map_req_v[700]));
	MUX21X1 U701(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[5]) ,.Q(int_map_req_v[701]));
	MUX21X1 U702(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[5]) ,.Q(int_map_req_v[702]));
	MUX21X1 U703(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[0]) ,.Q(int_map_req_v[703]));
	MUX21X1 U704(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[0]) ,.Q(int_map_req_v[704]));
	MUX21X1 U705(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[0]) ,.Q(int_map_req_v[705]));
	MUX21X1 U706(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[0]) ,.Q(int_map_req_v[706]));
	MUX21X1 U707(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[0]) ,.Q(int_map_req_v[707]));
	MUX21X1 U708(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[0]) ,.Q(int_map_req_v[708]));
	MUX21X1 U709(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[0]) ,.Q(int_map_req_v[709]));
	MUX21X1 U710(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[0]) ,.Q(int_map_req_v[710]));
	MUX21X1 U711(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[0]) ,.Q(int_map_req_v[711]));
	MUX21X1 U712(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[0]) ,.Q(int_map_req_v[712]));
	MUX21X1 U713(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[0]) ,.Q(int_map_req_v[713]));
	MUX21X1 U714(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[0]) ,.Q(int_map_req_v[714]));
	MUX21X1 U715(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[0]) ,.Q(int_map_req_v[715]));
	MUX21X1 U716(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[0]) ,.Q(int_map_req_v[716]));
	MUX21X1 U717(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[0]) ,.Q(int_map_req_v[717]));
	MUX21X1 U718(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[0]) ,.Q(int_map_req_v[718]));
	MUX21X1 U719(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[0]) ,.Q(int_map_req_v[719]));
	MUX21X1 U720(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[0]) ,.Q(int_map_req_v[720]));
	MUX21X1 U721(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[0]) ,.Q(int_map_req_v[721]));
	MUX21X1 U722(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[0]) ,.Q(int_map_req_v[722]));
	MUX21X1 U723(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[0]) ,.Q(int_map_req_v[723]));
	MUX21X1 U724(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[0]) ,.Q(int_map_req_v[724]));
	MUX21X1 U725(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[0]) ,.Q(int_map_req_v[725]));
	MUX21X1 U726(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[0]) ,.Q(int_map_req_v[726]));
	MUX21X1 U727(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[0]) ,.Q(int_map_req_v[727]));
	MUX21X1 U728(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[0]) ,.Q(int_map_req_v[728]));
	MUX21X1 U729(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[0]) ,.Q(int_map_req_v[729]));
	MUX21X1 U730(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[0]) ,.Q(int_map_req_v[730]));
	MUX21X1 U731(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[0]) ,.Q(int_map_req_v[731]));
	MUX21X1 U732(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[0]) ,.Q(int_map_req_v[732]));
	MUX21X1 U733(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[0]) ,.Q(int_map_req_v[733]));
	MUX21X1 U734(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[0]) ,.Q(int_map_req_v[734]));
	MUX21X1 U735(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[0]) ,.Q(int_map_req_v[735]));
	MUX21X1 U736(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[0]) ,.Q(int_map_req_v[736]));
	MUX21X1 U737(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[0]) ,.Q(int_map_req_v[737]));
	MUX21X1 U738(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[0]) ,.Q(int_map_req_v[738]));
	MUX21X1 U739(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[0]) ,.Q(int_map_req_v[739]));
	MUX21X1 U33(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[19]), .S(int_route_v[0]) ,.Q(int_resp_v[0]));
	MUX21X1 U34(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[20]), .S(int_route_v[0]) ,.Q(int_resp_v[1]));
	MUX21X1 U35(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[18]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));
	MUX21X1 U36(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[19]), .S(int_route_v[5]) ,.Q(int_resp_v[2]));
	MUX21X1 U37(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[17]), .S(int_route_v[10]) ,.Q(int_resp_v[2]));
	MUX21X1 U38(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[18]), .S(int_route_v[10]) ,.Q(int_resp_v[3]));
	MUX21X1 U39(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[16]), .S(int_route_v[15]) ,.Q(int_resp_v[3]));
	MUX21X1 U40(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[17]), .S(int_route_v[15]) ,.Q(int_resp_v[4]));
