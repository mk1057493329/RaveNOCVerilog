module router_ravenoc (clk,arst,north_send,north_recv,south_send,south_recv,west_send,west_recv,east_send,east_recv,local_send,local_recv);

	input clk;
	input arst;
	input north_send;
	input west_recv;
	input east_send;
	input east_recv;
	input north_recv;
	input south_send;
	input south_recv;
	input west_send;
	input local_send;
	input local_recv;
	
	wire south_recv_resp,south_recv_req,south_send_resp,south_send_req,west_recv_resp,west_recv_req,west_send_resp,west_send_req,north_recv_resp,north_recv_req,north_send_resp,north_send_req,east_recv_resp,east_recv_req,east_send_resp,east_send_req,local_recv_resp,local_recv_req,local_send_resp,local_send_req;
	wire [194:0] int_req_v;
	wire [4:0] int_resp_v;
	wire [24:0] int_route_v;
	wire [739:0] int_map_req_v;
	wire [19:0] int_map_resp_v;
	wire [194:0] ext_req_v_i;
	wire [4:0] ext_resp_v_o;
	wire [194:0] ext_req_v_o;
	wire [4:0] ext_resp_v_i;
	wire [11:0] valid_from_im_output_module;
	wire [11:0] grant_im_output_module;
	wire [2:0] tail_flit_im_output_module;
	wire [1:0] vc_ch_act_out_output_module;
	wire req_out_output_module,xnor1resu1_output_module,xnor2resu1_output_module,and1resu1_output_module,xor1resu1_output_module,and2resu1_output_module,head_flit_output_module_32_not_output_module,and3resu1_output_module,nor23resu1_output_module,nor23resu2_output_module,and4resu1_output_module,and5resu1_output_module,or12resu12_output_module,nor23resu3_output_module,and6resu1_output_module,nand1resu_output_module,and8resu1_output_module,norfinresu1_output_module,and9resu1_output_module,and10resu1_output_module,and11resu1_output_module;
	wire [33:0] head_flit_output_module;
	wire [1:0] _sv2v_jump_output_module;
	wire [31:0] in_mod_output_module;
	wire [31:0] vc_channel_output_module;
	wire [1:0] _sv2v_jump_output_module_1;
	wire [31:0] i_output_module;
    wire [1:0] mask_ff_rr_arbiter, next_mask_rr_arbiter, mask_req_rr_arbiter, _sv2v_jump_rr_rr_arbiter, i_rr_arbiter, j_rr_arbiter, raw_grant_rr_arbiter, masked_grant_rr_arbiter, temp_mask_ff_rr_arbiter, _sv2v_jump_high_prior_arbiter1, i_high_prior_arbiter1, _sv2v_jump_high_prior_arbiter2, i_high_prior_arbiter2, mask_ff_rr_arbiter1, next_mask_rr_arbiter1, mask_req_rr_arbiter1, _sv2v_jump_rr_rr_arbiter1, i_rr_arbiter1, j_rr_arbiter1, raw_grant_rr_arbiter1, masked_grant_rr_arbiter1, temp_mask_ff_rr_arbiter11, _sv2v_jump_high_prior_arbiter11, i_high_prior_arbiter11, _sv2v_jump_high_prior_arbiter21, i_high_prior_arbiter21,mask_ff_rr_arbiter2,next_mask_rr_arbiter2,mask_req_rr_arbiter2,_sv2v_jump_rr_rr_arbiter2,i_rr_arbiter2,j_rr_arbiter2,raw_grant_rr_arbiter2,masked_grant_rr_arbiter2,temp_mask_ff_rr_arbiter22,_sv2v_jump_high_prior_arbiter12,i_high_prior_arbiter12,_sv2v_jump_high_prior_arbiter22,i_high_prior_arbiter22;

    wire xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter,xnor1res_rr_arbiter,firstif_rr_arbiter,secondif_rr_arbiter,thirdif_rr_arbiter,fourthif_rr_arbiter,not_i_rr_arbiter,arst_value_rr_arbiter,xnores_high_prior_arbiter1,i_0_not_high_prior_arbiter1,nandres_high_prior_arbiter1,xnores_high_prior_arbiter2,i_0_not_high_prior_arbiter2,nandres_high_prior_arbiter2,xnor0res_rr_arbiter1,xnor1res_rr_arbiter1,firstif_rr_arbiter1,secondif_rr_arbiter1,thirdif_rr_arbiter1,fourthif_rr_arbiter1,not_i_rr_arbiter11,arst_value_rr_arbiter1,xnores_high_prior_arbiter11,i_0_not_high_prior_arbiter11,nandres_high_prior_arbiter11,xnores_high_prior_arbiter22,i_0_not_high_prior_arbiter22,nandres_high_prior_arbiter22,xnor0res_rr_arbiter2,xnor1res_rr_arbiter2,firstif_rr_arbiter2,secondif_rr_arbiter2,thirdif_rr_arbiter2,fourthif_rr_arbiter2,not_i_rr_arbiter22,arst_value_rr_arbiter2,xnores_high_prior_arbiter12,i_0_not_high_prior_arbiter12,nandres_high_prior_arbiter12;

    wire [11:0] valid_from_im_output_module1;
    wire [11:0] grant_im_output_module1;
    wire [2:0] tail_flit_im_output_module1;
    wire [1:0] vc_ch_act_out_output_module1;
    wire req_out_output_module1,xnor1resu1_output_module1,xnor2resu1_output_module1,and1resu1_output_module1,xor1resu1_output_module1,and2resu1_output_module1,head_flit_output_module1_32_not_output_module1,and3resu1_output_module1,nor23resu1_output_module1,nor23resu2_output_module1,and4resu1_output_module1,and5resu1_output_module1,or12resu12_output_module1,nor23resu3_output_module1,and6resu1_output_module1,nand1resu_output_module1,and8resu1_output_module1,norfinresu1_output_module1,and9resu1_output_module1,and10resu1_output_module1,and11resu1_output_module1;
    wire [33:0] head_flit_output_module1;
    wire [1:0] _sv2v_jump_output_module1;
    wire [31:0] in_mod_output_module1;
    wire [31:0] vc_channel_output_module1;
    wire [1:0] _sv2v_jump_output_module1_1;
    wire [31:0] i_output_module1;
    wire [1:0] mask_ff_rr_arbiter11, next_mask_rr_arbiter11, mask_req_rr_arbiter11, _sv2v_jump_rr_rr_arbiter11, i_rr_arbiter11, j_rr_arbiter11, raw_grant_rr_arbiter11, masked_grant_rr_arbiter11, temp_mask_ff_rr_arbiter1111, _sv2v_jump_high_prior_arbiter111, i_high_prior_arbiter111, _sv2v_jump_high_prior_arbiter211, i_high_prior_arbiter211, mask_ff_rr_arbiter111, next_mask_rr_arbiter111, mask_req_rr_arbiter111, _sv2v_jump_rr_rr_arbiter111, i_rr_arbiter111, j_rr_arbiter111, raw_grant_rr_arbiter111, masked_grant_rr_arbiter111, temp_mask_ff_rr_arbiter111111, _sv2v_jump_high_prior_arbiter1111, i_high_prior_arbiter1111, _sv2v_jump_high_prior_arbiter2111, i_high_prior_arbiter2111,mask_ff_rr_arbiter112,next_mask_rr_arbiter112,mask_req_rr_arbiter112,_sv2v_jump_rr_rr_arbiter112,i_rr_arbiter112,j_rr_arbiter112,raw_grant_rr_arbiter112,masked_grant_rr_arbiter112,temp_mask_ff_rr_arbiter111122,_sv2v_jump_high_prior_arbiter1112,i_high_prior_arbiter1112,_sv2v_jump_high_prior_arbiter2112,i_high_prior_arbiter2112;

    wire xnores_high_prior_arbiter2111,i_0_not_high_prior_arbiter2111,nandres_high_prior_arbiter2111,xnor0res_rr_arbiter11,xnor1res_rr_arbiter11,firstif_rr_arbiter11,secondif_rr_arbiter11,thirdif_rr_arbiter11,fourthif_rr_arbiter11,not_i_rr_arbiter1111,arst_value_rr_arbiter11,xnores_high_prior_arbiter111,i_0_not_high_prior_arbiter111,nandres_high_prior_arbiter111,xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter111,xnor1res_rr_arbiter111,firstif_rr_arbiter111,secondif_rr_arbiter111,thirdif_rr_arbiter111,fourthif_rr_arbiter111,not_i_rr_arbiter111111,arst_value_rr_arbiter111,xnores_high_prior_arbiter1111,i_0_not_high_prior_arbiter1111,nandres_high_prior_arbiter1111,xnores_high_prior_arbiter212,i_0_not_high_prior_arbiter212,nandres_high_prior_arbiter212,xnor0res_rr_arbiter112,xnor1res_rr_arbiter112,firstif_rr_arbiter112,secondif_rr_arbiter112,thirdif_rr_arbiter112,fourthif_rr_arbiter112,not_i_rr_arbiter111122,arst_value_rr_arbiter112,xnores_high_prior_arbiter1112,i_0_not_high_prior_arbiter1112,nandres_high_prior_arbiter1112;

    wire [11:0] valid_from_im_output_module2;
    wire [11:0] grant_im_output_module2;
    wire [2:0] tail_flit_im_output_module2;
    wire [1:0] vc_ch_act_out_output_module2;
    wire req_out_output_module2,xnor1resu1_output_module2,xnor2resu1_output_module2,and1resu1_output_module2,xor1resu1_output_module2,and2resu1_output_module2,head_flit_output_module2_32_not_output_module2,and3resu1_output_module2,nor23resu1_output_module2,nor23resu2_output_module2,and4resu1_output_module2,and5resu1_output_module2,or12resu12_output_module2,nor23resu3_output_module2,and6resu1_output_module2,nand1resu_output_module2,and8resu1_output_module2,norfinresu1_output_module2,and9resu1_output_module2,and10resu1_output_module2,and11resu1_output_module2;
    wire [33:0] head_flit_output_module2;
    wire [1:0] _sv2v_jump_output_module2;
    wire [31:0] in_mod_output_module2;
    wire [31:0] vc_channel_output_module2;
    wire [1:0] _sv2v_jump_output_module2_1;
    wire [31:0] i_output_module2;
    wire [1:0] mask_ff_rr_arbiter22, next_mask_rr_arbiter22, mask_req_rr_arbiter22, _sv2v_jump_rr_rr_arbiter22, i_rr_arbiter22, j_rr_arbiter22, raw_grant_rr_arbiter22, masked_grant_rr_arbiter22, temp_mask_ff_rr_arbiter2222, _sv2v_jump_high_prior_arbiter122, i_high_prior_arbiter122, _sv2v_jump_high_prior_arbiter222, i_high_prior_arbiter222, mask_ff_rr_arbiter221, next_mask_rr_arbiter221, mask_req_rr_arbiter221, _sv2v_jump_rr_rr_arbiter221, i_rr_arbiter221, j_rr_arbiter221, raw_grant_rr_arbiter221, masked_grant_rr_arbiter221, temp_mask_ff_rr_arbiter222211, _sv2v_jump_high_prior_arbiter1221, i_high_prior_arbiter1221, _sv2v_jump_high_prior_arbiter2221, i_high_prior_arbiter2221,mask_ff_rr_arbiter222,next_mask_rr_arbiter222,mask_req_rr_arbiter222,_sv2v_jump_rr_rr_arbiter222,i_rr_arbiter222,j_rr_arbiter222,raw_grant_rr_arbiter222,masked_grant_rr_arbiter222,temp_mask_ff_rr_arbiter222222,_sv2v_jump_high_prior_arbiter1222,i_high_prior_arbiter1222,_sv2v_jump_high_prior_arbiter2222,i_high_prior_arbiter2222;

    wire xnores_high_prior_arbiter22212,i_0_not_high_prior_arbiter22212,nandres_high_prior_arbiter22212,xnor0res_rr_arbiter22,xnor1res_rr_arbiter22,firstif_rr_arbiter22,secondif_rr_arbiter22,thirdif_rr_arbiter22,fourthif_rr_arbiter22,not_i_rr_arbiter2222,arst_value_rr_arbiter22,xnores_high_prior_arbiter122,i_0_not_high_prior_arbiter122,nandres_high_prior_arbiter122,xnores_high_prior_arbiter222,i_0_not_high_prior_arbiter222,nandres_high_prior_arbiter222,xnor0res_rr_arbiter221,xnor1res_rr_arbiter221,firstif_rr_arbiter221,secondif_rr_arbiter221,thirdif_rr_arbiter221,fourthif_rr_arbiter221,not_i_rr_arbiter222211,arst_value_rr_arbiter221,xnores_high_prior_arbiter1221,i_0_not_high_prior_arbiter1221,nandres_high_prior_arbiter1221,xnores_high_prior_arbiter2222,i_0_not_high_prior_arbiter2222,nandres_high_prior_arbiter2222,xnor0res_rr_arbiter222,xnor1res_rr_arbiter222,firstif_rr_arbiter222,secondif_rr_arbiter222,thirdif_rr_arbiter222,fourthif_rr_arbiter222,not_i_rr_arbiter222222,arst_value_rr_arbiter222,xnores_high_prior_arbiter1222,i_0_not_high_prior_arbiter1222,nandres_high_prior_arbiter1222;


    wire [11:0] valid_from_im_output_module3;
    wire [11:0] grant_im_output_module3;
    wire [2:0] tail_flit_im_output_module3;
    wire [1:0] vc_ch_act_out_output_module3;
    wire req_out_output_module3,xnor1resu1_output_module3,xnor2resu1_output_module3,and1resu1_output_module3,xor1resu1_output_module3,and2resu1_output_module3,head_flit_output_module3_32_not_output_module3,and3resu1_output_module3,nor23resu1_output_module3,nor23resu2_output_module3,and4resu1_output_module3,and5resu1_output_module3,or12resu12_output_module3,nor23resu3_output_module3,and6resu1_output_module3,nand1resu_output_module3,and8resu1_output_module3,norfinresu1_output_module3,and9resu1_output_module3,and10resu1_output_module3,and11resu1_output_module3;
    wire [33:0] head_flit_output_module3;
    wire [1:0] _sv2v_jump_output_module3;
    wire [31:0] in_mod_output_module3;
    wire [31:0] vc_channel_output_module3;
    wire [1:0] _sv2v_jump_output_module3_1;
    wire [31:0] i_output_module3;
    wire [1:0] mask_ff_rr_arbiter3, next_mask_rr_arbiter3, mask_req_rr_arbiter3, _sv2v_jump_rr_rr_arbiter3, i_rr_arbiter3, j_rr_arbiter3, raw_grant_rr_arbiter3, masked_grant_rr_arbiter3, temp_mask_ff_rr_arbiter33, _sv2v_jump_high_prior_arbiter13, i_high_prior_arbiter13, _sv2v_jump_high_prior_arbiter23, i_high_prior_arbiter23, mask_ff_rr_arbiter31, next_mask_rr_arbiter31, mask_req_rr_arbiter31, _sv2v_jump_rr_rr_arbiter31, i_rr_arbiter31, j_rr_arbiter31, raw_grant_rr_arbiter31, masked_grant_rr_arbiter31, temp_mask_ff_rr_arbiter3311, _sv2v_jump_high_prior_arbiter131, i_high_prior_arbiter131, _sv2v_jump_high_prior_arbiter231, i_high_prior_arbiter231,mask_ff_rr_arbiter32,next_mask_rr_arbiter32,mask_req_rr_arbiter32,_sv2v_jump_rr_rr_arbiter32,i_rr_arbiter32,j_rr_arbiter32,raw_grant_rr_arbiter32,masked_grant_rr_arbiter32,temp_mask_ff_rr_arbiter3322,_sv2v_jump_high_prior_arbiter132,i_high_prior_arbiter132,_sv2v_jump_high_prior_arbiter232,i_high_prior_arbiter232;

    wire xnores_high_prior_arbiter2313,i_0_not_high_prior_arbiter2313,nandres_high_prior_arbiter2313,xnor0res_rr_arbiter3,xnor1res_rr_arbiter3,firstif_rr_arbiter3,secondif_rr_arbiter3,thirdif_rr_arbiter3,fourthif_rr_arbiter3,not_i_rr_arbiter33,arst_value_rr_arbiter3,xnores_high_prior_arbiter13,i_0_not_high_prior_arbiter13,nandres_high_prior_arbiter13,xnores_high_prior_arbiter23,i_0_not_high_prior_arbiter23,nandres_high_prior_arbiter23,xnor0res_rr_arbiter31,xnor1res_rr_arbiter31,firstif_rr_arbiter31,secondif_rr_arbiter31,thirdif_rr_arbiter31,fourthif_rr_arbiter31,not_i_rr_arbiter3311,arst_value_rr_arbiter31,xnores_high_prior_arbiter131,i_0_not_high_prior_arbiter131,nandres_high_prior_arbiter131,xnores_high_prior_arbiter232,i_0_not_high_prior_arbiter232,nandres_high_prior_arbiter232,xnor0res_rr_arbiter32,xnor1res_rr_arbiter32,firstif_rr_arbiter32,secondif_rr_arbiter32,thirdif_rr_arbiter32,fourthif_rr_arbiter32,not_i_rr_arbiter3322,arst_value_rr_arbiter32,xnores_high_prior_arbiter132,i_0_not_high_prior_arbiter132,nandres_high_prior_arbiter132;


    wire [11:0] valid_from_im_output_module4;
    wire [11:0] grant_im_output_module4;
    wire [2:0] tail_flit_im_output_module4;
    wire [1:0] vc_ch_act_out_output_module4;
    wire req_out_output_module4,xnor1resu1_output_module4,xnor2resu1_output_module4,and1resu1_output_module4,xor1resu1_output_module4,and2resu1_output_module4,head_flit_output_module4_32_not_output_module4,and3resu1_output_module4,nor23resu1_output_module4,nor23resu2_output_module4,and4resu1_output_module4,and5resu1_output_module4,or12resu12_output_module4,nor23resu3_output_module4,and6resu1_output_module4,nand1resu_output_module4,and8resu1_output_module4,norfinresu1_output_module4,and9resu1_output_module4,and10resu1_output_module4,and11resu1_output_module4;
    wire [33:0] head_flit_output_module4;
    wire [1:0] _sv2v_jump_output_module4;
    wire [31:0] in_mod_output_module4;
    wire [31:0] vc_channel_output_module4;
    wire [1:0] _sv2v_jump_output_module4_1;
    wire [31:0] i_output_module4;
    wire [1:0] mask_ff_rr_arbiter4, next_mask_rr_arbiter4, mask_req_rr_arbiter4, _sv2v_jump_rr_rr_arbiter4, i_rr_arbiter4, j_rr_arbiter4, raw_grant_rr_arbiter4, masked_grant_rr_arbiter4, temp_mask_ff_rr_arbiter44, _sv2v_jump_high_prior_arbiter14, i_high_prior_arbiter14, _sv2v_jump_high_prior_arbiter24, i_high_prior_arbiter24, mask_ff_rr_arbiter41, next_mask_rr_arbiter41, mask_req_rr_arbiter41, _sv2v_jump_rr_rr_arbiter41, i_rr_arbiter41, j_rr_arbiter41, raw_grant_rr_arbiter41, masked_grant_rr_arbiter41, temp_mask_ff_rr_arbiter4411, _sv2v_jump_high_prior_arbiter141, i_high_prior_arbiter141, _sv2v_jump_high_prior_arbiter241, i_high_prior_arbiter241,mask_ff_rr_arbiter42,next_mask_rr_arbiter42,mask_req_rr_arbiter42,_sv2v_jump_rr_rr_arbiter42,i_rr_arbiter42,j_rr_arbiter42,raw_grant_rr_arbiter42,masked_grant_rr_arbiter42,temp_mask_ff_rr_arbiter4422,_sv2v_jump_high_prior_arbiter142,i_high_prior_arbiter142,_sv2v_jump_high_prior_arbiter242,i_high_prior_arbiter242;

    wire xnores_high_prior_arbiter2414,i_0_not_high_prior_arbiter2414,nandres_high_prior_arbiter2414,xnor0res_rr_arbiter4,xnor1res_rr_arbiter4,firstif_rr_arbiter4,secondif_rr_arbiter4,thirdif_rr_arbiter4,fourthif_rr_arbiter4,not_i_rr_arbiter44,arst_value_rr_arbiter4,xnores_high_prior_arbiter14,i_0_not_high_prior_arbiter14,nandres_high_prior_arbiter14,xnores_high_prior_arbiter24,i_0_not_high_prior_arbiter24,nandres_high_prior_arbiter24,xnor0res_rr_arbiter41,xnor1res_rr_arbiter41,firstif_rr_arbiter41,secondif_rr_arbiter41,thirdif_rr_arbiter41,fourthif_rr_arbiter41,not_i_rr_arbiter4411,arst_value_rr_arbiter41,xnores_high_prior_arbiter141,i_0_not_high_prior_arbiter141,nandres_high_prior_arbiter141,xnores_high_prior_arbiter242,i_0_not_high_prior_arbiter242,nandres_high_prior_arbiter242,xnor0res_rr_arbiter42,xnor1res_rr_arbiter42,firstif_rr_arbiter42,secondif_rr_arbiter42,thirdif_rr_arbiter42,fourthif_rr_arbiter42,not_i_rr_arbiter4422,arst_value_rr_arbiter42,xnores_high_prior_arbiter142,i_0_not_high_prior_arbiter142,nandres_high_prior_arbiter142;

   	wire [8:0] routing_table_ff_input_router;
	wire [2:0] next_rt_input_router;
	wire [33:0] flit_input_router;
	wire new_rt_input_router,new_rt_input_routernot,norres_1_input_router,norres_2_input_router,norres_3_input_router,andfinres_input_router,and2result_input_router,norres_4_input_router,invres1_input_router,invres2_input_router,and3result_input_router,and4result_input_router,and5result_input_router,norres_5_input_router,and6result_input_router,and7result_input_router,and8result_input_router,and9result_input_router,and10result_input_router,and11result_input_router,orres1_input_router,orres2_input_router,orres3_input_router,finand1_input_router,finand2_input_router,finand3_input_router,nextrt2not_input_router,secondAndc_input_router,norres_5_input_router_2,and62result_input_router,and7result_input_router2,orres1_input_router2,finand1_input_router2,finand2_input_router2,and8result_input_router2,orres2_input_router2,and9result_input_router2,orres3_input_router2,finand3_input_router2,and11result_input_router2,nextrt2not_input_router,and10result_input_router2,arst_valuenot_input_router,finand3_input_router22;
    
    wire [8:0] routing_table_ff_input_router1;
    wire [2:0] next_rt_input_router1;
    wire [33:0] flit_input_router1;
    wire new_rt_input_router1,new_rt_input_router1not,norres_1_input_router1,norres_2_input_router1,norres_3_input_router1,andfinres_input_router1,and2result_input_router1,norres_4_input_router1,invres1_input_router1,invres2_input_router1,and3result_input_router1,and4result_input_router1,and5result_input_router1,norres_5_input_router1,and6result_input_router1,and7result_input_router1,and8result_input_router1,and9result_input_router1,and10result_input_router1,and11result_input_router1,orres1_input_router1,orres2_input_router1,orres3_input_router1,finand1_input_router1,finand2_input_router1,finand3_input_router1,nextrt2not_input_router11,secondAndc_input_router1,norres_5_input_router1_2,and62result_input_router1,and7result_input_router12,orres1_input_router12,finand1_input_router12,finand2_input_router12,and8result_input_router12,orres2_input_router12,and9result_input_router12,orres3_input_router12,finand3_input_router12,and11result_input_router12,nextrt2not_input_router11,and10result_input_router12,arst_valuenot_input_router1,finand3_input_router122;


    wire [8:0] routing_table_ff_input_router2;
    wire [2:0] next_rt_input_router2;
    wire [33:0] flit_input_router2;
    wire new_rt_input_router2,new_rt_input_router2not,norres_1_input_router2,norres_2_input_router2,norres_3_input_router2,andfinres_input_router2,and2result_input_router2,norres_4_input_router2,invres1_input_router2,invres2_input_router2,and3result_input_router2,and4result_input_router2,and5result_input_router2,norres_5_input_router2,and6result_input_router2,and7result_input_router22,and8result_input_router22,and9result_input_router22,and10result_input_router22,and11result_input_router22,orres1_input_router22,orres2_input_router22,orres3_input_router22,finand1_input_router22,finand2_input_router22,finand3_input_router222,nextrt2not_input_router22,secondAndc_input_router2,norres_5_input_router2_2,and62result_input_router2,and7result_input_router222,orres1_input_router222,finand1_input_router222,finand2_input_router222,and8result_input_router222,orres2_input_router222,and9result_input_router222,orres3_input_router222,finand3_input_router2222,and11result_input_router222,nextrt2not_input_router22,and10result_input_router222,arst_valuenot_input_router2,finand3_input_router22222;


    wire [8:0] routing_table_ff_input_router3;
    wire [2:0] next_rt_input_router3;
    wire [33:0] flit_input_router3;
    wire new_rt_input_router3,new_rt_input_router3not,norres_1_input_router3,norres_2_input_router3,norres_3_input_router3,andfinres_input_router3,and2result_input_router3,norres_4_input_router3,invres1_input_router3,invres2_input_router3,and3result_input_router3,and4result_input_router3,and5result_input_router3,norres_5_input_router3,and6result_input_router3,and7result_input_router3,and8result_input_router3,and9result_input_router3,and10result_input_router3,and11result_input_router3,orres1_input_router3,orres2_input_router3,orres3_input_router3,finand1_input_router3,finand2_input_router3,finand3_input_router3,nextrt2not_input_router33,secondAndc_input_router3,norres_5_input_router3_2,and62result_input_router3,and7result_input_router32,orres1_input_router32,finand1_input_router32,finand2_input_router32,and8result_input_router32,orres2_input_router32,and9result_input_router32,orres3_input_router32,finand3_input_router32,and11result_input_router32,nextrt2not_input_router33,and10result_input_router32,arst_valuenot_input_router3,finand3_input_router322;


    wire [8:0] routing_table_ff_input_router4;
    wire [2:0] next_rt_input_router4;
    wire [33:0] flit_input_router4;
    wire new_rt_input_router4,new_rt_input_router4not,norres_1_input_router4,norres_2_input_router4,norres_3_input_router4,andfinres_input_router4,and2result_input_router4,norres_4_input_router4,invres1_input_router4,invres2_input_router4,and3result_input_router4,and4result_input_router4,and5result_input_router4,norres_5_input_router4,and6result_input_router4,and7result_input_router4,and8result_input_router4,and9result_input_router4,and10result_input_router4,and11result_input_router4,orres1_input_router4,orres2_input_router4,orres3_input_router4,finand1_input_router4,finand2_input_router4,finand3_input_router4,nextrt2not_input_router44,secondAndc_input_router4,norres_5_input_router4_2,and62result_input_router4,and7result_input_router42,orres1_input_router42,finand1_input_router42,finand2_input_router42,and8result_input_router42,orres2_input_router42,and9result_input_router42,orres3_input_router42,finand3_input_router42,and11result_input_router42,nextrt2not_input_router44,and10result_input_router42,arst_valuenot_input_router4,finand3_input_router422;

	wire [110:0] from_input_req_in_jump_input_datapathput_datapath;
	wire [2:0] from_input_resp_input_datapath;
	wire [110:0] to_output_req_in_jump_input_datapathput_datapath;
	wire [2:0] to_output_resp_input_datapath;
	wire [1:0] vc_ch_act_in_input_datapath;
	wire [1:0] vc_ch_act_out_input_datapath;
	wire [2:0] i_input_datapath;
	wire [2:0] j_input_datapath;
	wire [0:1] _sv2v_jump_input_datapath;

	wire req_in_jump_input_datapath,req_out_jump_input_datapath,xnor1resu_input_datapath,xnor2resu_input_datapath,and1resu_input_datapath,cond1line_input_datapath,req_in_jump_input_datapath_not,and2resu_input_datapath,xor1resu_input_datapath,nand1resu_input_datapath,xnor23resu_input_datapath,and4resu_input_datapath,write_flit_vc_buffer,norres_vc_buffer_vc_buffer,full_vc_buffer,empty_vc_buffer,error_vc_buffer,read_flit_vc_buffer,locked_by_route_ff_vc_buffer,next_locked_vc_buffer,orres_vc_buffer,or1res_vc_buffer,or2res_vc_buffer,finres1_vc_buffer,andres1_vc_buffer,full_vc_buffer_not,locked_by_route_ff_vc_buffer_not,thirdand_vc_buffer,u1temp_fifomodule,u2temp_fifomodule,u4temp_fifomodule,full_vc_buffer_not_fifomodule,u7temp_fifomodule,u9temp_fifomodule,u10carry_fifomodule,u11carry_fifomodule,empty_vc_buffer_not_fifomodule,u13temp_fifomodule,u14temp_fifomodule,u15carry_fifomodule,u16carry_fifomodule,u17res_fifomodule,u18res_fifomodule,write_ptr_ff_fifomodule_0_not,write_ptr_ff_fifomodule_1_not,b0wire_fifomodule,b1wire_fifomodule,u23temp_fifomodule_not_fifomodule,u23temp_fifomodule,boutb_fifomodule,bouta_fifomodule,boutmain_fifomodule,arst_value_fifomodule,write_flit1_vc_buffer1,norres_vc_buffer1_vc_buffer1,full_vc_buffer1,empty_vc_buffer1,error_vc_buffer1,read_flit1_vc_buffer1,locked_by_route_ff_vc_buffer1,next_locked_vc_buffer1,orres_vc_buffer1,or1res_vc_buffer1,or2res_vc_buffer1,finres1_vc_buffer1,andres1_vc_buffer1,full_vc_buffer1_not1,locked_by_route_ff_vc_buffer1_not1,thirdand_vc_buffer1,u1temp_fifomodule1,u2temp_fifomodule1,u4temp_fifomodule1,full_vc_buffer1_not1_fifomodule1,u7temp_fifomodule1,u9temp_fifomodule1,u10carry_fifomodule1,u11carry_fifomodule1,empty_vc_buffer1_not_fifomodule1,u13temp_fifomodule1,u14temp_fifomodule1,u15carry_fifomodule1,u16carry_fifomodule1,u17res_fifomodule1,u18res_fifomodule1,write_ptr_ff_fifomodule1_0_not1,write_ptr_ff_fifomodule1_1_not1,b0wire_fifomodule1,b1wire_fifomodule1,u23temp_fifomodule1_not_fifomodule1,u23temp_fifomodule1,boutb_fifomodule1,bouta_fifomodule1,boutmain_fifomodule1,arst_value_fifomodule1,write_flit2_vc_buffer2,norres_vc_buffer2_vc_buffer2,full_vc_buffer2,empty_vc_buffer2,error_vc_buffer2,read_flit2_vc_buffer2,locked_by_route_ff_vc_buffer2,next_locked_vc_buffer2,orres_vc_buffer2,or1res_vc_buffer2,or2res_vc_buffer2,finres1_vc_buffer2,andres1_vc_buffer2,full_vc_buffer2_not2,locked_by_route_ff_vc_buffer2_not2,thirdand_vc_buffer2,u1temp_fifomodule2,u2temp_fifomodule2,u4temp_fifomodule2,full_vc_buffer2_not2_fifomodule2,u7temp_fifomodule2,u9temp_fifomodule2,u10carry_fifomodule2,u11carry_fifomodule2,empty_vc_buffer2_not_fifomodule2,u13temp_fifomodule2,u14temp_fifomodule2,u15carry_fifomodule2,u16carry_fifomodule2,u17res_fifomodule2,u18res_fifomodule2,write_ptr_ff_fifomodule2_0_not2,write_ptr_ff_fifomodule2_1_not2,b0wire_fifomodule2,b1wire_fifomodule2,u23temp_fifomodule2_not_fifomodule2,u23temp_fifomodule2,boutb_fifomodule2,bouta_fifomodule2,boutmain_fifomodule2,arst_value_fifomodule2;
	wire [33:0] flit,flit1,flit2;
	wire [15:0] fifo_ff_fifomodule,fifo_ff_fifomodule1,fifo_ff_fifomodule2;
	wire [1:0] write_ptr_ff_fifomodule,read_ptr_ff_fifomodule,next_write_ptr_fifomodule,next_read_ptr_fifomodule,fifo_ocup_fifomodule,write_ptr_ff_fifomodule1,read_ptr_ff_fifomodule1,next_write_ptr_fifomodule1,next_read_ptr_fifomodule1,fifo_ocup_fifomodule1,write_ptr_ff_fifomodule2,read_ptr_ff_fifomodule2,next_write_ptr_fifomodule2,next_read_ptr_fifomodule2,fifo_ocup_fifomodule2;

	wire [110:0] from_input_req_in_jump_input_datapath1put_datapath1;
	wire [2:0] from_input_resp_input_datapath1;
	wire [110:0] to_output_req_in_jump_input_datapath1put_datapath1;
	wire [2:0] to_output_resp_input_datapath1;
	wire [1:0] vc_ch_act_in_input_datapath1;
	wire [1:0] vc_ch_act_out_input_datapath1;
	wire [2:0] i_input_datapath1;
	wire [2:0] j_input_datapath1;
	wire [0:1] _sv2v_jump_input_datapath1;

	wire req_in_jump_input_datapath1,req_out_jump_input_datapath1,xnor1resu_input_datapath1,xnor2resu_input_datapath1,and1resu_input_datapath1,cond1line_input_datapath1,req_in_jump_input_datapath1_not,and2resu_input_datapath1,xor1resu_input_datapath1,nand1resu_input_datapath11,xnor23resu_input_datapath1,and4resu_input_datapath1,write_flit11_vc_buffer1,norres_vc_buffer11_vc_buffer11,full_vc_buffer11,empty_vc_buffer11,error_vc_buffer11,read_flit11_vc_buffer1,locked_by_route_ff_vc_buffer11,next_locked_vc_buffer11,orres_vc_buffer11,or1res_vc_buffer11,or2res_vc_buffer11,finres1_vc_buffer11,andres1_vc_buffer11,full_vc_buffer11_not,locked_by_route_ff_vc_buffer11_not,thirdand_vc_buffer11,u1temp_fifomodule11,u2temp_fifomodule11,u4temp_fifomodule11,full_vc_buffer11_not_fifomodule,u7temp_fifomodule11,u9temp_fifomodule11,u10carry_fifomodule11,u11carry_fifomodule11,empty_vc_buffer11_not_fifomodule,u13temp_fifomodule11,u14temp_fifomodule11,u15carry_fifomodule11,u16carry_fifomodule11,u17res_fifomodule11,u18res_fifomodule11,write_ptr_ff_fifomodule11_0_not1,write_ptr_ff_fifomodule11_1_not1,b0wire_fifomodule11,b1wire_fifomodule11,u23temp_fifomodule11_not_fifomodule11,u23temp_fifomodule11,boutb_fifomodule11,bouta_fifomodule11,boutmain_fifomodule11,arst_value_fifomodule11,write_flit111_vc_buffer11,norres_vc_buffer111_vc_buffer1,full_vc_buffer111,empty_vc_buffer111,error_vc_buffer111,read_flit111_vc_buffer11,locked_by_route_ff_vc_buffer111,next_locked_vc_buffer111,orres_vc_buffer111,or1res_vc_buffer111,or2res_vc_buffer111,finres1_vc_buffer111,andres1_vc_buffer111,full_vc_buffer111_not1,locked_by_route_ff_vc_buffer111_not1,thirdand_vc_buffer111,u1temp_fifomodule111,u2temp_fifomodule111,u4temp_fifomodule111,full_vc_buffer111_not1_fifomodule1,u7temp_fifomodule111,u9temp_fifomodule111,u10carry_fifomodule111,u11carry_fifomodule111,empty_vc_buffer111_not_fifomodule1,u13temp_fifomodule111,u14temp_fifomodule111,u15carry_fifomodule111,u16carry_fifomodule111,u17res_fifomodule111,u18res_fifomodule111,write_ptr_ff_fifomodule111_0_not11,write_ptr_ff_fifomodule111_1_not11,b0wire_fifomodule111,b1wire_fifomodule111,u23temp_fifomodule111_not_fifomodule1,u23temp_fifomodule111,boutb_fifomodule111,bouta_fifomodule111,boutmain_fifomodule111,arst_value_fifomodule111,write_flit112_vc_buffer21,norres_vc_buffer112_vc_buffer2,full_vc_buffer112,empty_vc_buffer112,error_vc_buffer112,read_flit112_vc_buffer21,locked_by_route_ff_vc_buffer112,next_locked_vc_buffer112,orres_vc_buffer112,or1res_vc_buffer112,or2res_vc_buffer112,finres1_vc_buffer112,andres1_vc_buffer112,full_vc_buffer112_not2,locked_by_route_ff_vc_buffer112_not2,thirdand_vc_buffer112,u1temp_fifomodule112,u2temp_fifomodule112,u4temp_fifomodule112,full_vc_buffer112_not2_fifomodule2,u7temp_fifomodule112,u9temp_fifomodule112,u10carry_fifomodule112,u11carry_fifomodule112,empty_vc_buffer112_not_fifomodule2,u13temp_fifomodule112,u14temp_fifomodule112,u15carry_fifomodule112,u16carry_fifomodule112,u17res_fifomodule112,u18res_fifomodule112,write_ptr_ff_fifomodule112_0_not21,write_ptr_ff_fifomodule112_1_not21,b0wire_fifomodule112,b1wire_fifomodule112,u23temp_fifomodule112_not_fifomodule2,u23temp_fifomodule112,boutb_fifomodule112,bouta_fifomodule112,boutmain_fifomodule112,arst_value_fifomodule112;
	wire [33:0] flit11,flit111,flit112;
	wire [15:0] fifo_ff_fifomodule11,fifo_ff_fifomodule111,fifo_ff_fifomodule112;
	wire [1:0] write_ptr_ff_fifomodule11,read_ptr_ff_fifomodule11,next_write_ptr_fifomodule11,next_read_ptr_fifomodule11,fifo_ocup_fifomodule11,write_ptr_ff_fifomodule111,read_ptr_ff_fifomodule111,next_write_ptr_fifomodule111,next_read_ptr_fifomodule111,fifo_ocup_fifomodule111,write_ptr_ff_fifomodule112,read_ptr_ff_fifomodule112,next_write_ptr_fifomodule112,next_read_ptr_fifomodule112,fifo_ocup_fifomodule112;

	wire [110:0] from_input_req_in_jump_input_datapath2put_datapath2;
	wire [2:0] from_input_resp_input_datapath2;
	wire [110:0] to_output_req_in_jump_input_datapath2put_datapath2;
	wire [2:0] to_output_resp_input_datapath2;
	wire [1:0] vc_ch_act_in_input_datapath2;
	wire [1:0] vc_ch_act_out_input_datapath2;
	wire [2:0] i_input_datapath2;
	wire [2:0] j_input_datapath2;
	wire [0:1] _sv2v_jump_input_datapath2;

	wire req_in_jump_input_datapath2,req_out_jump_input_datapath2,xnor1resu_input_datapath2,xnor2resu_input_datapath2,and1resu_input_datapath2,cond1line_input_datapath2,req_in_jump_input_datapath2_not,and2resu_input_datapath2,xor1resu_input_datapath2,nand1resu_input_datapath22,xnor23resu_input_datapath2,and4resu_input_datapath2,write_flit22_vc_buffer2,norres_vc_buffer22_vc_buffer22,full_vc_buffer22,empty_vc_buffer22,error_vc_buffer22,read_flit22_vc_buffer2,locked_by_route_ff_vc_buffer22,next_locked_vc_buffer22,orres_vc_buffer22,or1res_vc_buffer22,or2res_vc_buffer22,finres1_vc_buffer22,andres1_vc_buffer22,full_vc_buffer22_not,locked_by_route_ff_vc_buffer22_not,thirdand_vc_buffer22,u1temp_fifomodule22,u2temp_fifomodule22,u4temp_fifomodule22,full_vc_buffer22_not_fifomodule,u7temp_fifomodule22,u9temp_fifomodule22,u10carry_fifomodule22,u11carry_fifomodule22,empty_vc_buffer22_not_fifomodule,u13temp_fifomodule22,u14temp_fifomodule22,u15carry_fifomodule22,u16carry_fifomodule22,u17res_fifomodule22,u18res_fifomodule22,write_ptr_ff_fifomodule22_0_not2,write_ptr_ff_fifomodule22_1_not2,b0wire_fifomodule22,b1wire_fifomodule22,u23temp_fifomodule22_not_fifomodule22,u23temp_fifomodule22,boutb_fifomodule22,bouta_fifomodule22,boutmain_fifomodule22,arst_value_fifomodule22,write_flit221_vc_buffer12,norres_vc_buffer221_vc_buffer1,full_vc_buffer221,empty_vc_buffer221,error_vc_buffer221,read_flit221_vc_buffer12,locked_by_route_ff_vc_buffer221,next_locked_vc_buffer221,orres_vc_buffer221,or1res_vc_buffer221,or2res_vc_buffer221,finres1_vc_buffer221,andres1_vc_buffer221,full_vc_buffer221_not1,locked_by_route_ff_vc_buffer221_not1,thirdand_vc_buffer221,u1temp_fifomodule221,u2temp_fifomodule221,u4temp_fifomodule221,full_vc_buffer221_not1_fifomodule1,u7temp_fifomodule221,u9temp_fifomodule221,u10carry_fifomodule221,u11carry_fifomodule221,empty_vc_buffer221_not_fifomodule1,u13temp_fifomodule221,u14temp_fifomodule221,u15carry_fifomodule221,u16carry_fifomodule221,u17res_fifomodule221,u18res_fifomodule221,write_ptr_ff_fifomodule221_0_not12,write_ptr_ff_fifomodule221_1_not12,b0wire_fifomodule221,b1wire_fifomodule221,u23temp_fifomodule221_not_fifomodule1,u23temp_fifomodule221,boutb_fifomodule221,bouta_fifomodule221,boutmain_fifomodule221,arst_value_fifomodule221,write_flit222_vc_buffer22,norres_vc_buffer222_vc_buffer2,full_vc_buffer222,empty_vc_buffer222,error_vc_buffer222,read_flit222_vc_buffer22,locked_by_route_ff_vc_buffer222,next_locked_vc_buffer222,orres_vc_buffer222,or1res_vc_buffer222,or2res_vc_buffer222,finres1_vc_buffer222,andres1_vc_buffer222,full_vc_buffer222_not2,locked_by_route_ff_vc_buffer222_not2,thirdand_vc_buffer222,u1temp_fifomodule222,u2temp_fifomodule222,u4temp_fifomodule222,full_vc_buffer222_not2_fifomodule2,u7temp_fifomodule222,u9temp_fifomodule222,u10carry_fifomodule222,u11carry_fifomodule222,empty_vc_buffer222_not_fifomodule2,u13temp_fifomodule222,u14temp_fifomodule222,u15carry_fifomodule222,u16carry_fifomodule222,u17res_fifomodule222,u18res_fifomodule222,write_ptr_ff_fifomodule222_0_not22,write_ptr_ff_fifomodule222_1_not22,b0wire_fifomodule222,b1wire_fifomodule222,u23temp_fifomodule222_not_fifomodule2,u23temp_fifomodule222,boutb_fifomodule222,bouta_fifomodule222,boutmain_fifomodule222,arst_value_fifomodule222;
	wire [33:0] flit22,flit221,flit222;
	wire [15:0] fifo_ff_fifomodule22,fifo_ff_fifomodule221,fifo_ff_fifomodule222;
	wire [1:0] write_ptr_ff_fifomodule22,read_ptr_ff_fifomodule22,next_write_ptr_fifomodule22,next_read_ptr_fifomodule22,fifo_ocup_fifomodule22,write_ptr_ff_fifomodule221,read_ptr_ff_fifomodule221,next_write_ptr_fifomodule221,next_read_ptr_fifomodule221,fifo_ocup_fifomodule221,write_ptr_ff_fifomodule222,read_ptr_ff_fifomodule222,next_write_ptr_fifomodule222,next_read_ptr_fifomodule222,fifo_ocup_fifomodule222;

	wire [110:0] from_input_req_in_jump_input_datapath3put_datapath3;
	wire [2:0] from_input_resp_input_datapath3;
	wire [110:0] to_output_req_in_jump_input_datapath3put_datapath3;
	wire [2:0] to_output_resp_input_datapath3;
	wire [1:0] vc_ch_act_in_input_datapath3;
	wire [1:0] vc_ch_act_out_input_datapath3;
	wire [2:0] i_input_datapath3;
	wire [2:0] j_input_datapath3;
	wire [0:1] _sv2v_jump_input_datapath3;

	wire req_in_jump_input_datapath3,req_out_jump_input_datapath3,xnor1resu_input_datapath3,xnor2resu_input_datapath3,and1resu_input_datapath3,cond1line_input_datapath3,req_in_jump_input_datapath3_not,and2resu_input_datapath3,xor1resu_input_datapath3,nand1resu_input_datapath33,xnor23resu_input_datapath3,and4resu_input_datapath3,write_flit3_vc_buffer3,norres_vc_buffer3_vc_buffer3,full_vc_buffer3,empty_vc_buffer3,error_vc_buffer3,read_flit3_vc_buffer3,locked_by_route_ff_vc_buffer3,next_locked_vc_buffer3,orres_vc_buffer3,or1res_vc_buffer3,or2res_vc_buffer3,finres1_vc_buffer3,andres1_vc_buffer3,full_vc_buffer3_not,locked_by_route_ff_vc_buffer3_not,thirdand_vc_buffer3,u1temp_fifomodule3,u2temp_fifomodule3,u4temp_fifomodule3,full_vc_buffer3_not_fifomodule,u7temp_fifomodule3,u9temp_fifomodule3,u10carry_fifomodule3,u11carry_fifomodule3,empty_vc_buffer3_not_fifomodule,u13temp_fifomodule3,u14temp_fifomodule3,u15carry_fifomodule3,u16carry_fifomodule3,u17res_fifomodule3,u18res_fifomodule3,write_ptr_ff_fifomodule3_0_not3,write_ptr_ff_fifomodule3_1_not3,b0wire_fifomodule3,b1wire_fifomodule3,u23temp_fifomodule3_not_fifomodule3,u23temp_fifomodule3,boutb_fifomodule3,bouta_fifomodule3,boutmain_fifomodule3,arst_value_fifomodule3,write_flit31_vc_buffer13,norres_vc_buffer31_vc_buffer1,full_vc_buffer31,empty_vc_buffer31,error_vc_buffer31,read_flit31_vc_buffer13,locked_by_route_ff_vc_buffer31,next_locked_vc_buffer31,orres_vc_buffer31,or1res_vc_buffer31,or2res_vc_buffer31,finres1_vc_buffer31,andres1_vc_buffer31,full_vc_buffer31_not1,locked_by_route_ff_vc_buffer31_not1,thirdand_vc_buffer31,u1temp_fifomodule31,u2temp_fifomodule31,u4temp_fifomodule31,full_vc_buffer31_not1_fifomodule1,u7temp_fifomodule31,u9temp_fifomodule31,u10carry_fifomodule31,u11carry_fifomodule31,empty_vc_buffer31_not_fifomodule1,u13temp_fifomodule31,u14temp_fifomodule31,u15carry_fifomodule31,u16carry_fifomodule31,u17res_fifomodule31,u18res_fifomodule31,write_ptr_ff_fifomodule31_0_not13,write_ptr_ff_fifomodule31_1_not13,b0wire_fifomodule31,b1wire_fifomodule31,u23temp_fifomodule31_not_fifomodule1,u23temp_fifomodule31,boutb_fifomodule31,bouta_fifomodule31,boutmain_fifomodule31,arst_value_fifomodule31,write_flit32_vc_buffer23,norres_vc_buffer32_vc_buffer2,full_vc_buffer32,empty_vc_buffer32,error_vc_buffer32,read_flit32_vc_buffer23,locked_by_route_ff_vc_buffer32,next_locked_vc_buffer32,orres_vc_buffer32,or1res_vc_buffer32,or2res_vc_buffer32,finres1_vc_buffer32,andres1_vc_buffer32,full_vc_buffer32_not2,locked_by_route_ff_vc_buffer32_not2,thirdand_vc_buffer32,u1temp_fifomodule32,u2temp_fifomodule32,u4temp_fifomodule32,full_vc_buffer32_not2_fifomodule2,u7temp_fifomodule32,u9temp_fifomodule32,u10carry_fifomodule32,u11carry_fifomodule32,empty_vc_buffer32_not_fifomodule2,u13temp_fifomodule32,u14temp_fifomodule32,u15carry_fifomodule32,u16carry_fifomodule32,u17res_fifomodule32,u18res_fifomodule32,write_ptr_ff_fifomodule32_0_not23,write_ptr_ff_fifomodule32_1_not23,b0wire_fifomodule32,b1wire_fifomodule32,u23temp_fifomodule32_not_fifomodule2,u23temp_fifomodule32,boutb_fifomodule32,bouta_fifomodule32,boutmain_fifomodule32,arst_value_fifomodule32;
	wire [33:0] flit3,flit31,flit32;
	wire [15:0] fifo_ff_fifomodule3,fifo_ff_fifomodule31,fifo_ff_fifomodule32;
	wire [1:0] write_ptr_ff_fifomodule3,read_ptr_ff_fifomodule3,next_write_ptr_fifomodule3,next_read_ptr_fifomodule3,fifo_ocup_fifomodule3,write_ptr_ff_fifomodule31,read_ptr_ff_fifomodule31,next_write_ptr_fifomodule31,next_read_ptr_fifomodule31,fifo_ocup_fifomodule31,write_ptr_ff_fifomodule32,read_ptr_ff_fifomodule32,next_write_ptr_fifomodule32,next_read_ptr_fifomodule32,fifo_ocup_fifomodule32;


	wire [110:0] from_input_req_in_jump_input_datapath4put_datapath4;
	wire [2:0] from_input_resp_input_datapath4;
	wire [110:0] to_output_req_in_jump_input_datapath4put_datapath4;
	wire [2:0] to_output_resp_input_datapath4;
	wire [1:0] vc_ch_act_in_input_datapath4;
	wire [1:0] vc_ch_act_out_input_datapath4;
	wire [2:0] i_input_datapath4;
	wire [2:0] j_input_datapath4;
	wire [0:1] _sv2v_jump_input_datapath4;

	wire req_in_jump_input_datapath4,req_out_jump_input_datapath4,xnor1resu_input_datapath4,xnor2resu_input_datapath4,and1resu_input_datapath4,cond1line_input_datapath4,req_in_jump_input_datapath4_not,and2resu_input_datapath4,xor1resu_input_datapath4,nand1resu_input_datapath44,xnor23resu_input_datapath4,and4resu_input_datapath4,write_flit4_vc_buffer4,norres_vc_buffer4_vc_buffer4,full_vc_buffer4,empty_vc_buffer4,error_vc_buffer4,read_flit4_vc_buffer4,locked_by_route_ff_vc_buffer4,next_locked_vc_buffer4,orres_vc_buffer4,or1res_vc_buffer4,or2res_vc_buffer4,finres1_vc_buffer4,andres1_vc_buffer4,full_vc_buffer4_not,locked_by_route_ff_vc_buffer4_not,thirdand_vc_buffer4,u1temp_fifomodule4,u2temp_fifomodule4,u4temp_fifomodule4,full_vc_buffer4_not_fifomodule,u7temp_fifomodule4,u9temp_fifomodule4,u10carry_fifomodule4,u11carry_fifomodule4,empty_vc_buffer4_not_fifomodule,u13temp_fifomodule4,u14temp_fifomodule4,u15carry_fifomodule4,u16carry_fifomodule4,u17res_fifomodule4,u18res_fifomodule4,write_ptr_ff_fifomodule4_0_not4,write_ptr_ff_fifomodule4_1_not4,b0wire_fifomodule4,b1wire_fifomodule4,u23temp_fifomodule4_not_fifomodule4,u23temp_fifomodule4,boutb_fifomodule4,bouta_fifomodule4,boutmain_fifomodule4,arst_value_fifomodule4,write_flit41_vc_buffer14,norres_vc_buffer41_vc_buffer1,full_vc_buffer41,empty_vc_buffer41,error_vc_buffer41,read_flit41_vc_buffer14,locked_by_route_ff_vc_buffer41,next_locked_vc_buffer41,orres_vc_buffer41,or1res_vc_buffer41,or2res_vc_buffer41,finres1_vc_buffer41,andres1_vc_buffer41,full_vc_buffer41_not1,locked_by_route_ff_vc_buffer41_not1,thirdand_vc_buffer41,u1temp_fifomodule41,u2temp_fifomodule41,u4temp_fifomodule41,full_vc_buffer41_not1_fifomodule1,u7temp_fifomodule41,u9temp_fifomodule41,u10carry_fifomodule41,u11carry_fifomodule41,empty_vc_buffer41_not_fifomodule1,u13temp_fifomodule41,u14temp_fifomodule41,u15carry_fifomodule41,u16carry_fifomodule41,u17res_fifomodule41,u18res_fifomodule41,write_ptr_ff_fifomodule41_0_not14,write_ptr_ff_fifomodule41_1_not14,b0wire_fifomodule41,b1wire_fifomodule41,u23temp_fifomodule41_not_fifomodule1,u23temp_fifomodule41,boutb_fifomodule41,bouta_fifomodule41,boutmain_fifomodule41,arst_value_fifomodule41,write_flit42_vc_buffer24,norres_vc_buffer42_vc_buffer2,full_vc_buffer42,empty_vc_buffer42,error_vc_buffer42,read_flit42_vc_buffer24,locked_by_route_ff_vc_buffer42,next_locked_vc_buffer42,orres_vc_buffer42,or1res_vc_buffer42,or2res_vc_buffer42,finres1_vc_buffer42,andres1_vc_buffer42,full_vc_buffer42_not2,locked_by_route_ff_vc_buffer42_not2,thirdand_vc_buffer42,u1temp_fifomodule42,u2temp_fifomodule42,u4temp_fifomodule42,full_vc_buffer42_not2_fifomodule2,u7temp_fifomodule42,u9temp_fifomodule42,u10carry_fifomodule42,u11carry_fifomodule42,empty_vc_buffer42_not_fifomodule2,u13temp_fifomodule42,u14temp_fifomodule42,u15carry_fifomodule42,u16carry_fifomodule42,u17res_fifomodule42,u18res_fifomodule42,write_ptr_ff_fifomodule42_0_not24,write_ptr_ff_fifomodule42_1_not24,b0wire_fifomodule42,b1wire_fifomodule42,u23temp_fifomodule42_not_fifomodule2,u23temp_fifomodule42,boutb_fifomodule42,bouta_fifomodule42,boutmain_fifomodule42,arst_value_fifomodule42;
	wire [33:0] flit4,flit41,flit42;
	wire [15:0] fifo_ff_fifomodule4,fifo_ff_fifomodule41,fifo_ff_fifomodule42;
	wire [1:0] write_ptr_ff_fifomodule4,read_ptr_ff_fifomodule4,next_write_ptr_fifomodule4,next_read_ptr_fifomodule4,fifo_ocup_fifomodule4,write_ptr_ff_fifomodule41,read_ptr_ff_fifomodule41,next_write_ptr_fifomodule41,next_read_ptr_fifomodule41,fifo_ocup_fifomodule41,write_ptr_ff_fifomodule42,read_ptr_ff_fifomodule42,next_write_ptr_fifomodule42,next_read_ptr_fifomodule42,fifo_ocup_fifomodule42;



//input router
    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router[2]) );
    BUFX1 U3(.A(flit_input_router_req_i[3]), .Y(flit_input_router[3]));
	BUFX1 U4(.A(flit_input_router_req_i[4]), .Y(flit_input_router[4]));
	BUFX1 U5(.A(flit_input_router_req_i[5]), .Y(flit_input_router[5]));
	BUFX1 U6(.A(flit_input_router_req_i[6]), .Y(flit_input_router[6]));
	BUFX1 U7(.A(flit_input_router_req_i[7]), .Y(flit_input_router[7]));
	BUFX1 U8(.A(flit_input_router_req_i[8]), .Y(flit_input_router[8]));
	BUFX1 U9(.A(flit_input_router_req_i[9]), .Y(flit_input_router[9]));
	BUFX1 U10(.A(flit_input_router_req_i[10]), .Y(flit_input_router[10]));
	BUFX1 U11(.A(flit_input_router_req_i[11]), .Y(flit_input_router[11]));
	BUFX1 U12(.A(flit_input_router_req_i[12]), .Y(flit_input_router[12]));
	BUFX1 U13(.A(flit_input_router_req_i[13]), .Y(flit_input_router[13]));
	BUFX1 U14(.A(flit_input_router_req_i[14]), .Y(flit_input_router[14]));
	BUFX1 U15(.A(flit_input_router_req_i[15]), .Y(flit_input_router[15]));
	BUFX1 U16(.A(flit_input_router_req_i[16]), .Y(flit_input_router[16]));
	BUFX1 U17(.A(flit_input_router_req_i[17]), .Y(flit_input_router[17]));
	BUFX1 U18(.A(flit_input_router_req_i[18]), .Y(flit_input_router[18]));
	BUFX1 U19(.A(flit_input_router_req_i[19]), .Y(flit_input_router[19]));
	BUFX1 U20(.A(flit_input_router_req_i[20]), .Y(flit_input_router[20]));
	BUFX1 U21(.A(flit_input_router_req_i[21]), .Y(flit_input_router[21]));
	BUFX1 U22(.A(flit_input_router_req_i[22]), .Y(flit_input_router[22]));
	BUFX1 U23(.A(flit_input_router_req_i[23]), .Y(flit_input_router[23]));
	BUFX1 U24(.A(flit_input_router_req_i[24]), .Y(flit_input_router[24]));
	BUFX1 U25(.A(flit_input_router_req_i[25]), .Y(flit_input_router[25]));
	BUFX1 U26(.A(flit_input_router_req_i[26]), .Y(flit_input_router[26]));
	BUFX1 U27(.A(flit_input_router_req_i[27]), .Y(flit_input_router[27]));
	BUFX1 U28(.A(flit_input_router_req_i[28]), .Y(flit_input_router[28]));
	BUFX1 U29(.A(flit_input_router_req_i[29]), .Y(flit_input_router[29]));
	BUFX1 U30(.A(flit_input_router_req_i[30]), .Y(flit_input_router[30]));
	BUFX1 U31(.A(flit_input_router_req_i[31]), .Y(flit_input_router[31]));
	BUFX1 U32(.A(flit_input_router_req_i[32]), .Y(flit_input_router[32]));
	BUFX1 U33(.A(flit_input_router_req_i[33]), .Y(flit_input_router[33]));
	BUFX1 U34(.A(flit_input_router_req_i[34]), .Y(flit_input_router[34]));
	BUFX1 U35(.A(flit_input_router_req_i[35]), .Y(flit_input_router[35]));
	BUFX1 U36(.A(flit_input_router_req_i[36]), .Y(flit_input_router[36]));

    NOR2X1 U37 ( .IN1(flit_input_router[33]), .IN2(flit_input_router[32]), .QN(norres_1_input_router) );
    AND2X1 U38 ( .IN1(flit_input_router_req_i[0]), .IN2(norres_1_input_router), .Q(new_rt_input_router) );

    NOR2X1 U37 ( .IN1(flit_input_router[31]), .IN2(1'b0), .QN(norres_2_input_router) );
    NOR2X1 U37 ( .IN1(flit_input_router[30]), .IN2(1'b0), .QN(norres_3_input_router) );
    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(norres_3_input_router), .Q(andfinres_input_router) );
    MUX21X1 U38 (.IN1(next_rt_input_router[0]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router[1]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router[2]), .IN2(1'b1), .S(andfinres_input_router), .Q(next_rt_input_router[2]);
    INVX1 U41 ( .A(andfinres_input_router), .Y(invres1_input_router) );


    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(invres1_input_router), .Q(and2result_input_router) );
    MUX21X1 U38 (.IN1(next_rt_input_router[0]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router[1]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router[2]), .IN2(1'b0), .S(and2result_input_router), .Q(next_rt_input_router[2]);
    INVX1 U41 ( .A(and2result_input_router), .Y(invres2_input_router) );

    AND3X1 U37 ( .IN1(new_rt_input_router), .IN2(invres1_input_router), .IN3(invres2_input_router), .Q(and3result_input_router) );
    AND2X1 U38 ( .IN1(flit_input_router[31]), .IN2(1'b1), .Q(and4result_input_router) );
    AND2X1 U38 ( .IN1(and4result_input_router), .IN2(and3result_input_router), .Q(and5result_input_router) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[2]);

   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][0]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][1]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][2]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][3]));
   	BUFX1 U35(.A(1'sb0), .Y(int_route_v[4:0][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(norres_5_input_router) );
    AND2X1 U38 ( .IN1(norres_5_input_router), .IN2(new_rt_input_router), .Q(and6result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and6result_input_router), .Q(int_route_v[4:0][4]);

    NOR2X1 U38 ( .IN1(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(and7result_input_router) );
    AND2X1 U19 ( .IN1(and7result_input_router), .IN2(next_rt_input_router[0]), .Y(orres1_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres1_input_router), .Q(finand1_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router), .Q(int_route_v[4:0][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[2]), .Q(and8result_input_router) );
    AND2X1 U19 ( .IN1(and8result_input_router), .IN2(next_rt_input_router[1]), .Y(orres2_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres2_input_router), .Q(finand2_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router), .Q(int_route_v[4:0][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and9result_input_router) );
    AND2X1 U19 ( .IN1(and9result_input_router), .IN2(next_rt_input_router[2]), .Y(orres3_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(orres3_input_router), .Q(finand3_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router), .Q(int_route_v[4:0][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and10result_input_router) );
    INVX1 U41 ( .A(next_rt_input_router[2]), .Y(nextrt2not_input_router) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router), .Q(and11result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    INVX1 U41 ( .A(new_rt_input_router), .Y(new_rt_input_routernot) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(flit_input_router_req_i[0]), .Q(secondAndc_input_router) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(norres_5_input_router_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router_2), .IN2(newsecondAndc_input_router_rt), .Q(and62result_input_router) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and62result_input_router), .Q(int_route_v[4:0][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(and7result_input_router2) );
    AND2X1 U19 ( .IN1(and7result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .Y(orres1_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres1_input_router2), .Q(finand1_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router2), .Q(int_route_v[4:0][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Q(and8result_input_router2) );
    AND2X1 U19 ( .IN1(and8result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Y(orres2_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres2_input_router), .Q(finand2_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router2), .Q(int_route_v[4:0][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and9result_input_router2) );
    AND2X1 U19 ( .IN1(and9result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(orres3_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_routernot), .IN2(orres3_input_router2), .Q(finand3_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router2), .Q(int_route_v[4:0][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and10result_input_router2) );
    INVX1 U41 ( .A(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(nextrt2not_input_router) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router2), .IN3(new_rt_input_routernot), .Q(and11result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router) );
    AND2X1 U38 ( .IN1(new_rt_input_router), .IN2(arst_valuenot_input_router), .Q(finand3_input_router22) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(next_rt_input_router[0]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(next_rt_input_router[1]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .IN2(next_rt_input_router[2]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]);    

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router1[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router1[2]) );
    BUFX1 U3(.A(flit_input_router1_req_i[3]), .Y(flit_input_router1[3]));
    BUFX1 U4(.A(flit_input_router1_req_i[4]), .Y(flit_input_router1[4]));
    BUFX1 U5(.A(flit_input_router1_req_i[5]), .Y(flit_input_router1[5]));
    BUFX1 U6(.A(flit_input_router1_req_i[6]), .Y(flit_input_router1[6]));
    BUFX1 U7(.A(flit_input_router1_req_i[7]), .Y(flit_input_router1[7]));
    BUFX1 U8(.A(flit_input_router1_req_i[8]), .Y(flit_input_router1[8]));
    BUFX1 U9(.A(flit_input_router1_req_i[9]), .Y(flit_input_router1[9]));
    BUFX1 U10(.A(flit_input_router1_req_i[10]), .Y(flit_input_router1[10]));
    BUFX1 U11(.A(flit_input_router1_req_i[11]), .Y(flit_input_router1[11]));
    BUFX1 U12(.A(flit_input_router1_req_i[12]), .Y(flit_input_router1[12]));
    BUFX1 U13(.A(flit_input_router1_req_i[13]), .Y(flit_input_router1[13]));
    BUFX1 U14(.A(flit_input_router1_req_i[14]), .Y(flit_input_router1[14]));
    BUFX1 U15(.A(flit_input_router1_req_i[15]), .Y(flit_input_router1[15]));
    BUFX1 U16(.A(flit_input_router1_req_i[16]), .Y(flit_input_router1[16]));
    BUFX1 U17(.A(flit_input_router1_req_i[17]), .Y(flit_input_router1[17]));
    BUFX1 U18(.A(flit_input_router1_req_i[18]), .Y(flit_input_router1[18]));
    BUFX1 U19(.A(flit_input_router1_req_i[19]), .Y(flit_input_router1[19]));
    BUFX1 U20(.A(flit_input_router1_req_i[20]), .Y(flit_input_router1[20]));
    BUFX1 U21(.A(flit_input_router1_req_i[21]), .Y(flit_input_router1[21]));
    BUFX1 U22(.A(flit_input_router1_req_i[22]), .Y(flit_input_router1[22]));
    BUFX1 U23(.A(flit_input_router1_req_i[23]), .Y(flit_input_router1[23]));
    BUFX1 U24(.A(flit_input_router1_req_i[24]), .Y(flit_input_router1[24]));
    BUFX1 U25(.A(flit_input_router1_req_i[25]), .Y(flit_input_router1[25]));
    BUFX1 U26(.A(flit_input_router1_req_i[26]), .Y(flit_input_router1[26]));
    BUFX1 U27(.A(flit_input_router1_req_i[27]), .Y(flit_input_router1[27]));
    BUFX1 U28(.A(flit_input_router1_req_i[28]), .Y(flit_input_router1[28]));
    BUFX1 U29(.A(flit_input_router1_req_i[29]), .Y(flit_input_router1[29]));
    BUFX1 U30(.A(flit_input_router1_req_i[30]), .Y(flit_input_router1[30]));
    BUFX1 U31(.A(flit_input_router1_req_i[31]), .Y(flit_input_router1[31]));
    BUFX1 U32(.A(flit_input_router1_req_i[32]), .Y(flit_input_router1[32]));
    BUFX1 U33(.A(flit_input_router1_req_i[33]), .Y(flit_input_router1[33]));
    BUFX1 U34(.A(flit_input_router1_req_i[34]), .Y(flit_input_router1[34]));
    BUFX1 U35(.A(flit_input_router1_req_i[35]), .Y(flit_input_router1[35]));
    BUFX1 U36(.A(flit_input_router1_req_i[36]), .Y(flit_input_router1[36]));

    NOR2X1 U37 ( .IN1(flit_input_router1[33]), .IN2(flit_input_router1[32]), .QN(norres_1_input_router1) );
    AND2X1 U38 ( .IN1(flit_input_router1_req_i[0]), .IN2(norres_1_input_router1), .Q(new_rt_input_router1) );

    NOR2X1 U37 ( .IN1(flit_input_router1[31]), .IN2(1'b0), .QN(norres_2_input_router1) );
    NOR2X1 U37 ( .IN1(flit_input_router1[30]), .IN2(1'b0), .QN(norres_3_input_router1) );
    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(norres_3_input_router1), .Q(andfinres_input_router1) );
    MUX21X1 U38 (.IN1(next_rt_input_router1[0]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[1]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[2]), .IN2(1'b1), .S(andfinres_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U41 ( .A(andfinres_input_router1), .Y(invres1_input_router1) );


    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(invres1_input_router1), .Q(and2result_input_router1) );
    MUX21X1 U38 (.IN1(next_rt_input_router1[0]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[1]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router1[2]), .IN2(1'b0), .S(and2result_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U41 ( .A(and2result_input_router1), .Y(invres2_input_router1) );

    AND3X1 U37 ( .IN1(new_rt_input_router1), .IN2(invres1_input_router1), .IN3(invres2_input_router1), .Q(and3result_input_router1) );
    AND2X1 U38 ( .IN1(flit_input_router1[31]), .IN2(1'b1), .Q(and4result_input_router1) );
    AND2X1 U38 ( .IN1(and4result_input_router1), .IN2(and3result_input_router1), .Q(and5result_input_router1) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[9:5][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(norres_5_input_router1) );
    AND2X1 U38 ( .IN1(norres_5_input_router1), .IN2(new_rt_input_router1), .Q(and6result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and6result_input_router1), .Q(int_route_v[9:5][4]);

    NOR2X1 U38 ( .IN1(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(and7result_input_router1) );
    AND2X1 U19 ( .IN1(and7result_input_router1), .IN2(next_rt_input_router1[0]), .Y(orres1_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres1_input_router1), .Q(finand1_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router1), .Q(int_route_v[9:5][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[2]), .Q(and8result_input_router1) );
    AND2X1 U19 ( .IN1(and8result_input_router1), .IN2(next_rt_input_router1[1]), .Y(orres2_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres2_input_router1), .Q(finand2_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router1), .Q(int_route_v[9:5][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and9result_input_router1) );
    AND2X1 U19 ( .IN1(and9result_input_router1), .IN2(next_rt_input_router1[2]), .Y(orres3_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(orres3_input_router1), .Q(finand3_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router1), .Q(int_route_v[9:5][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and10result_input_router1) );
    INVX1 U41 ( .A(next_rt_input_router1[2]), .Y(nextrt2not_input_router11) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router1), .Q(and11result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    INVX1 U41 ( .A(new_rt_input_router1), .Y(new_rt_input_router1not) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(flit_input_router1_req_i[0]), .Q(secondAndc_input_router1) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(norres_5_input_router1_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router1_2), .IN2(newsecondAndc_input_router1_rt), .Q(and62result_input_router1) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and62result_input_router1), .Q(int_route_v[9:5][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(and7result_input_router12) );
    AND2X1 U19 ( .IN1(and7result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .Y(orres1_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres1_input_router12), .Q(finand1_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router12), .Q(int_route_v[9:5][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Q(and8result_input_router12) );
    AND2X1 U19 ( .IN1(and8result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Y(orres2_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres2_input_router1), .Q(finand2_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router12), .Q(int_route_v[9:5][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and9result_input_router12) );
    AND2X1 U19 ( .IN1(and9result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(orres3_input_router12) );
    AND2X1 U38 ( .IN1(new_rt_input_router1not), .IN2(orres3_input_router12), .Q(finand3_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router12), .Q(int_route_v[9:5][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and10result_input_router12) );
    INVX1 U41 ( .A(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(nextrt2not_input_router11) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router12), .IN3(new_rt_input_router1not), .Q(and11result_input_router12) );
    MUX21X1 U38 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router1) );
    AND2X1 U38 ( .IN1(new_rt_input_router1), .IN2(arst_valuenot_input_router1), .Q(finand3_input_router122) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(next_rt_input_router1[0]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(next_rt_input_router1[1]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .IN2(next_rt_input_router1[2]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]);


	BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router2[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router2[2]) );
    BUFX1 U3(.A(flit_input_router2_req_i[3]), .Y(flit_input_router2[3]));
    BUFX1 U4(.A(flit_input_router2_req_i[4]), .Y(flit_input_router2[4]));
    BUFX1 U5(.A(flit_input_router2_req_i[5]), .Y(flit_input_router2[5]));
    BUFX1 U6(.A(flit_input_router2_req_i[6]), .Y(flit_input_router2[6]));
    BUFX1 U7(.A(flit_input_router2_req_i[7]), .Y(flit_input_router2[7]));
    BUFX1 U8(.A(flit_input_router2_req_i[8]), .Y(flit_input_router2[8]));
    BUFX1 U9(.A(flit_input_router2_req_i[9]), .Y(flit_input_router2[9]));
    BUFX1 U10(.A(flit_input_router2_req_i[10]), .Y(flit_input_router2[10]));
    BUFX1 U11(.A(flit_input_router2_req_i[11]), .Y(flit_input_router2[11]));
    BUFX1 U12(.A(flit_input_router2_req_i[12]), .Y(flit_input_router2[12]));
    BUFX1 U13(.A(flit_input_router2_req_i[13]), .Y(flit_input_router2[13]));
    BUFX1 U14(.A(flit_input_router2_req_i[14]), .Y(flit_input_router2[14]));
    BUFX1 U15(.A(flit_input_router2_req_i[15]), .Y(flit_input_router2[15]));
    BUFX1 U16(.A(flit_input_router2_req_i[16]), .Y(flit_input_router2[16]));
    BUFX1 U17(.A(flit_input_router2_req_i[17]), .Y(flit_input_router2[17]));
    BUFX1 U18(.A(flit_input_router2_req_i[18]), .Y(flit_input_router2[18]));
    BUFX1 U19(.A(flit_input_router2_req_i[19]), .Y(flit_input_router2[19]));
    BUFX1 U20(.A(flit_input_router2_req_i[20]), .Y(flit_input_router2[20]));
    BUFX1 U21(.A(flit_input_router2_req_i[21]), .Y(flit_input_router2[21]));
    BUFX1 U22(.A(flit_input_router2_req_i[22]), .Y(flit_input_router2[22]));
    BUFX1 U23(.A(flit_input_router2_req_i[23]), .Y(flit_input_router2[23]));
    BUFX1 U24(.A(flit_input_router2_req_i[24]), .Y(flit_input_router2[24]));
    BUFX1 U25(.A(flit_input_router2_req_i[25]), .Y(flit_input_router2[25]));
    BUFX1 U26(.A(flit_input_router2_req_i[26]), .Y(flit_input_router2[26]));
    BUFX1 U27(.A(flit_input_router2_req_i[27]), .Y(flit_input_router2[27]));
    BUFX1 U28(.A(flit_input_router2_req_i[28]), .Y(flit_input_router2[28]));
    BUFX1 U29(.A(flit_input_router2_req_i[29]), .Y(flit_input_router2[29]));
    BUFX1 U30(.A(flit_input_router2_req_i[30]), .Y(flit_input_router2[30]));
    BUFX1 U31(.A(flit_input_router2_req_i[31]), .Y(flit_input_router2[31]));
    BUFX1 U32(.A(flit_input_router2_req_i[32]), .Y(flit_input_router2[32]));
    BUFX1 U33(.A(flit_input_router2_req_i[33]), .Y(flit_input_router2[33]));
    BUFX1 U34(.A(flit_input_router2_req_i[34]), .Y(flit_input_router2[34]));
    BUFX1 U35(.A(flit_input_router2_req_i[35]), .Y(flit_input_router2[35]));
    BUFX1 U36(.A(flit_input_router2_req_i[36]), .Y(flit_input_router2[36]));

    NOR2X1 U37 ( .IN1(flit_input_router2[33]), .IN2(flit_input_router2[32]), .QN(norres_1_input_router2) );
    AND2X1 U38 ( .IN1(flit_input_router2_req_i[0]), .IN2(norres_1_input_router2), .Q(new_rt_input_router2) );

    NOR2X1 U37 ( .IN1(flit_input_router2[31]), .IN2(1'b0), .QN(norres_2_input_router2) );
    NOR2X1 U37 ( .IN1(flit_input_router2[30]), .IN2(1'b0), .QN(norres_3_input_router2) );
    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(norres_3_input_router2), .Q(andfinres_input_router2) );
    MUX21X1 U38 (.IN1(next_rt_input_router2[0]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[1]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[2]), .IN2(1'b1), .S(andfinres_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U41 ( .A(andfinres_input_router2), .Y(invres1_input_router2) );


    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(invres1_input_router2), .Q(and2result_input_router2) );
    MUX21X1 U38 (.IN1(next_rt_input_router2[0]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[1]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router2[2]), .IN2(1'b0), .S(and2result_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U41 ( .A(and2result_input_router2), .Y(invres2_input_router2) );

    AND3X1 U37 ( .IN1(new_rt_input_router2), .IN2(invres1_input_router2), .IN3(invres2_input_router2), .Q(and3result_input_router2) );
    AND2X1 U38 ( .IN1(flit_input_router2[31]), .IN2(1'b1), .Q(and4result_input_router2) );
    AND2X1 U38 ( .IN1(and4result_input_router2), .IN2(and3result_input_router2), .Q(and5result_input_router2) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[14:10][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(norres_5_input_router2) );
    AND2X1 U38 ( .IN1(norres_5_input_router2), .IN2(new_rt_input_router2), .Q(and6result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and6result_input_router2), .Q(int_route_v[14:10][4]);

    NOR2X1 U38 ( .IN1(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(and7result_input_router22) );
    AND2X1 U19 ( .IN1(and7result_input_router22), .IN2(next_rt_input_router2[0]), .Y(orres1_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres1_input_router22), .Q(finand1_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router22), .Q(int_route_v[14:10][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[2]), .Q(and8result_input_router22) );
    AND2X1 U19 ( .IN1(and8result_input_router22), .IN2(next_rt_input_router2[1]), .Y(orres2_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres2_input_router22), .Q(finand2_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router22), .Q(int_route_v[14:10][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and9result_input_router22) );
    AND2X1 U19 ( .IN1(and9result_input_router22), .IN2(next_rt_input_router2[2]), .Y(orres3_input_router22) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(orres3_input_router22), .Q(finand3_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router222), .Q(int_route_v[14:10][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and10result_input_router22) );
    INVX1 U41 ( .A(next_rt_input_router2[2]), .Y(nextrt2not_input_router22) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router22), .Q(and11result_input_router22) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    INVX1 U41 ( .A(new_rt_input_router2), .Y(new_rt_input_router2not) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(flit_input_router2_req_i[0]), .Q(secondAndc_input_router2) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(norres_5_input_router2_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router2_2), .IN2(newsecondAndc_input_router2_rt), .Q(and62result_input_router2) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and62result_input_router2), .Q(int_route_v[14:10][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(and7result_input_router222) );
    AND2X1 U19 ( .IN1(and7result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .Y(orres1_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres1_input_router222), .Q(finand1_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router222), .Q(int_route_v[14:10][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Q(and8result_input_router222) );
    AND2X1 U19 ( .IN1(and8result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Y(orres2_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres2_input_router22), .Q(finand2_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router222), .Q(int_route_v[14:10][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and9result_input_router222) );
    AND2X1 U19 ( .IN1(and9result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(orres3_input_router222) );
    AND2X1 U38 ( .IN1(new_rt_input_router2not), .IN2(orres3_input_router222), .Q(finand3_input_router2222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router2222), .Q(int_route_v[14:10][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and10result_input_router222) );
    INVX1 U41 ( .A(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(nextrt2not_input_router22) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router222), .IN3(new_rt_input_router2not), .Q(and11result_input_router222) );
    MUX21X1 U38 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router2) );
    AND2X1 U38 ( .IN1(new_rt_input_router2), .IN2(arst_valuenot_input_router2), .Q(finand3_input_router22222) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(next_rt_input_router2[0]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(next_rt_input_router2[1]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .IN2(next_rt_input_router2[2]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]); 

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router3[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router3[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router3[2]) );
    BUFX1 U3(.A(flit_input_router3_req_i[3]), .Y(flit_input_router3[3]));
    BUFX1 U4(.A(flit_input_router3_req_i[4]), .Y(flit_input_router3[4]));
    BUFX1 U5(.A(flit_input_router3_req_i[5]), .Y(flit_input_router3[5]));
    BUFX1 U6(.A(flit_input_router3_req_i[6]), .Y(flit_input_router3[6]));
    BUFX1 U7(.A(flit_input_router3_req_i[7]), .Y(flit_input_router3[7]));
    BUFX1 U8(.A(flit_input_router3_req_i[8]), .Y(flit_input_router3[8]));
    BUFX1 U9(.A(flit_input_router3_req_i[9]), .Y(flit_input_router3[9]));
    BUFX1 U10(.A(flit_input_router3_req_i[10]), .Y(flit_input_router3[10]));
    BUFX1 U11(.A(flit_input_router3_req_i[11]), .Y(flit_input_router3[11]));
    BUFX1 U12(.A(flit_input_router3_req_i[12]), .Y(flit_input_router3[12]));
    BUFX1 U13(.A(flit_input_router3_req_i[13]), .Y(flit_input_router3[13]));
    BUFX1 U14(.A(flit_input_router3_req_i[14]), .Y(flit_input_router3[14]));
    BUFX1 U15(.A(flit_input_router3_req_i[15]), .Y(flit_input_router3[15]));
    BUFX1 U16(.A(flit_input_router3_req_i[16]), .Y(flit_input_router3[16]));
    BUFX1 U17(.A(flit_input_router3_req_i[17]), .Y(flit_input_router3[17]));
    BUFX1 U18(.A(flit_input_router3_req_i[18]), .Y(flit_input_router3[18]));
    BUFX1 U19(.A(flit_input_router3_req_i[19]), .Y(flit_input_router3[19]));
    BUFX1 U20(.A(flit_input_router3_req_i[20]), .Y(flit_input_router3[20]));
    BUFX1 U21(.A(flit_input_router3_req_i[21]), .Y(flit_input_router3[21]));
    BUFX1 U22(.A(flit_input_router3_req_i[22]), .Y(flit_input_router3[22]));
    BUFX1 U23(.A(flit_input_router3_req_i[23]), .Y(flit_input_router3[23]));
    BUFX1 U24(.A(flit_input_router3_req_i[24]), .Y(flit_input_router3[24]));
    BUFX1 U25(.A(flit_input_router3_req_i[25]), .Y(flit_input_router3[25]));
    BUFX1 U26(.A(flit_input_router3_req_i[26]), .Y(flit_input_router3[26]));
    BUFX1 U27(.A(flit_input_router3_req_i[27]), .Y(flit_input_router3[27]));
    BUFX1 U28(.A(flit_input_router3_req_i[28]), .Y(flit_input_router3[28]));
    BUFX1 U29(.A(flit_input_router3_req_i[29]), .Y(flit_input_router3[29]));
    BUFX1 U30(.A(flit_input_router3_req_i[30]), .Y(flit_input_router3[30]));
    BUFX1 U31(.A(flit_input_router3_req_i[31]), .Y(flit_input_router3[31]));
    BUFX1 U32(.A(flit_input_router3_req_i[32]), .Y(flit_input_router3[32]));
    BUFX1 U33(.A(flit_input_router3_req_i[33]), .Y(flit_input_router3[33]));
    BUFX1 U34(.A(flit_input_router3_req_i[34]), .Y(flit_input_router3[34]));
    BUFX1 U35(.A(flit_input_router3_req_i[35]), .Y(flit_input_router3[35]));
    BUFX1 U36(.A(flit_input_router3_req_i[36]), .Y(flit_input_router3[36]));

    NOR2X1 U37 ( .IN1(flit_input_router3[33]), .IN2(flit_input_router3[32]), .QN(norres_1_input_router3) );
    AND2X1 U38 ( .IN1(flit_input_router3_req_i[0]), .IN2(norres_1_input_router3), .Q(new_rt_input_router3) );

    NOR2X1 U37 ( .IN1(flit_input_router3[31]), .IN2(1'b0), .QN(norres_2_input_router3) );
    NOR2X1 U37 ( .IN1(flit_input_router3[30]), .IN2(1'b0), .QN(norres_3_input_router3) );
    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(norres_3_input_router3), .Q(andfinres_input_router3) );
    MUX21X1 U38 (.IN1(next_rt_input_router3[0]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[1]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[2]), .IN2(1'b1), .S(andfinres_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U41 ( .A(andfinres_input_router3), .Y(invres1_input_router3) );


    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(invres1_input_router3), .Q(and2result_input_router3) );
    MUX21X1 U38 (.IN1(next_rt_input_router3[0]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[1]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router3[2]), .IN2(1'b0), .S(and2result_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U41 ( .A(and2result_input_router3), .Y(invres2_input_router3) );

    AND3X1 U37 ( .IN1(new_rt_input_router3), .IN2(invres1_input_router3), .IN3(invres2_input_router3), .Q(and3result_input_router3) );
    AND2X1 U38 ( .IN1(flit_input_router3[31]), .IN2(1'b1), .Q(and4result_input_router3) );
    AND2X1 U38 ( .IN1(and4result_input_router3), .IN2(and3result_input_router3), .Q(and5result_input_router3) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[19:15][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(norres_5_input_router3) );
    AND2X1 U38 ( .IN1(norres_5_input_router3), .IN2(new_rt_input_router3), .Q(and6result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and6result_input_router3), .Q(int_route_v[19:15][4]);

    NOR2X1 U38 ( .IN1(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(and7result_input_router3) );
    AND2X1 U19 ( .IN1(and7result_input_router3), .IN2(next_rt_input_router3[0]), .Y(orres1_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres1_input_router3), .Q(finand1_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router3), .Q(int_route_v[19:15][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[2]), .Q(and8result_input_router3) );
    AND2X1 U19 ( .IN1(and8result_input_router3), .IN2(next_rt_input_router3[1]), .Y(orres2_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres2_input_router3), .Q(finand2_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router3), .Q(int_route_v[19:15][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and9result_input_router3) );
    AND2X1 U19 ( .IN1(and9result_input_router3), .IN2(next_rt_input_router3[2]), .Y(orres3_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(orres3_input_router3), .Q(finand3_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router3), .Q(int_route_v[19:15][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and10result_input_router3) );
    INVX1 U41 ( .A(next_rt_input_router3[2]), .Y(nextrt2not_input_router33) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router3), .Q(and11result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    INVX1 U41 ( .A(new_rt_input_router3), .Y(new_rt_input_router3not) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(flit_input_router3_req_i[0]), .Q(secondAndc_input_router3) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(norres_5_input_router3_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router3_2), .IN2(newsecondAndc_input_router3_rt), .Q(and62result_input_router3) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and62result_input_router3), .Q(int_route_v[19:15][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(and7result_input_router32) );
    AND2X1 U19 ( .IN1(and7result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .Y(orres1_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres1_input_router32), .Q(finand1_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router32), .Q(int_route_v[19:15][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Q(and8result_input_router32) );
    AND2X1 U19 ( .IN1(and8result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Y(orres2_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres2_input_router3), .Q(finand2_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router32), .Q(int_route_v[19:15][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and9result_input_router32) );
    AND2X1 U19 ( .IN1(and9result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(orres3_input_router32) );
    AND2X1 U38 ( .IN1(new_rt_input_router3not), .IN2(orres3_input_router32), .Q(finand3_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router32), .Q(int_route_v[19:15][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and10result_input_router32) );
    INVX1 U41 ( .A(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(nextrt2not_input_router33) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router32), .IN3(new_rt_input_router3not), .Q(and11result_input_router32) );
    MUX21X1 U38 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router3) );
    AND2X1 U38 ( .IN1(new_rt_input_router3), .IN2(arst_valuenot_input_router3), .Q(finand3_input_router322) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(next_rt_input_router3[0]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(next_rt_input_router3[1]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .IN2(next_rt_input_router3[2]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]);

    BUFX1 U00 ( .A(1'b0), .Y(next_rt_input_router4[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(next_rt_input_router4[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(next_rt_input_router4[2]) );
    BUFX1 U3(.A(flit_input_router4_req_i[3]), .Y(flit_input_router4[3]));
    BUFX1 U4(.A(flit_input_router4_req_i[4]), .Y(flit_input_router4[4]));
    BUFX1 U5(.A(flit_input_router4_req_i[5]), .Y(flit_input_router4[5]));
    BUFX1 U6(.A(flit_input_router4_req_i[6]), .Y(flit_input_router4[6]));
    BUFX1 U7(.A(flit_input_router4_req_i[7]), .Y(flit_input_router4[7]));
    BUFX1 U8(.A(flit_input_router4_req_i[8]), .Y(flit_input_router4[8]));
    BUFX1 U9(.A(flit_input_router4_req_i[9]), .Y(flit_input_router4[9]));
    BUFX1 U10(.A(flit_input_router4_req_i[10]), .Y(flit_input_router4[10]));
    BUFX1 U11(.A(flit_input_router4_req_i[11]), .Y(flit_input_router4[11]));
    BUFX1 U12(.A(flit_input_router4_req_i[12]), .Y(flit_input_router4[12]));
    BUFX1 U13(.A(flit_input_router4_req_i[13]), .Y(flit_input_router4[13]));
    BUFX1 U14(.A(flit_input_router4_req_i[14]), .Y(flit_input_router4[14]));
    BUFX1 U15(.A(flit_input_router4_req_i[15]), .Y(flit_input_router4[15]));
    BUFX1 U16(.A(flit_input_router4_req_i[16]), .Y(flit_input_router4[16]));
    BUFX1 U17(.A(flit_input_router4_req_i[17]), .Y(flit_input_router4[17]));
    BUFX1 U18(.A(flit_input_router4_req_i[18]), .Y(flit_input_router4[18]));
    BUFX1 U19(.A(flit_input_router4_req_i[19]), .Y(flit_input_router4[19]));
    BUFX1 U20(.A(flit_input_router4_req_i[20]), .Y(flit_input_router4[20]));
    BUFX1 U21(.A(flit_input_router4_req_i[21]), .Y(flit_input_router4[21]));
    BUFX1 U22(.A(flit_input_router4_req_i[22]), .Y(flit_input_router4[22]));
    BUFX1 U23(.A(flit_input_router4_req_i[23]), .Y(flit_input_router4[23]));
    BUFX1 U24(.A(flit_input_router4_req_i[24]), .Y(flit_input_router4[24]));
    BUFX1 U25(.A(flit_input_router4_req_i[25]), .Y(flit_input_router4[25]));
    BUFX1 U26(.A(flit_input_router4_req_i[26]), .Y(flit_input_router4[26]));
    BUFX1 U27(.A(flit_input_router4_req_i[27]), .Y(flit_input_router4[27]));
    BUFX1 U28(.A(flit_input_router4_req_i[28]), .Y(flit_input_router4[28]));
    BUFX1 U29(.A(flit_input_router4_req_i[29]), .Y(flit_input_router4[29]));
    BUFX1 U30(.A(flit_input_router4_req_i[30]), .Y(flit_input_router4[30]));
    BUFX1 U31(.A(flit_input_router4_req_i[31]), .Y(flit_input_router4[31]));
    BUFX1 U32(.A(flit_input_router4_req_i[32]), .Y(flit_input_router4[32]));
    BUFX1 U33(.A(flit_input_router4_req_i[33]), .Y(flit_input_router4[33]));
    BUFX1 U34(.A(flit_input_router4_req_i[34]), .Y(flit_input_router4[34]));
    BUFX1 U35(.A(flit_input_router4_req_i[35]), .Y(flit_input_router4[35]));
    BUFX1 U36(.A(flit_input_router4_req_i[36]), .Y(flit_input_router4[36]));

    NOR2X1 U37 ( .IN1(flit_input_router4[33]), .IN2(flit_input_router4[32]), .QN(norres_1_input_router4) );
    AND2X1 U38 ( .IN1(flit_input_router4_req_i[0]), .IN2(norres_1_input_router4), .Q(new_rt_input_router4) );

    NOR2X1 U37 ( .IN1(flit_input_router4[31]), .IN2(1'b0), .QN(norres_2_input_router4) );
    NOR2X1 U37 ( .IN1(flit_input_router4[30]), .IN2(1'b0), .QN(norres_3_input_router4) );
    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(norres_3_input_router4), .Q(andfinres_input_router4) );
    MUX21X1 U38 (.IN1(next_rt_input_router4[0]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[1]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[2]), .IN2(1'b1), .S(andfinres_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U41 ( .A(andfinres_input_router4), .Y(invres1_input_router4) );


    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(invres1_input_router4), .Q(and2result_input_router4) );
    MUX21X1 U38 (.IN1(next_rt_input_router4[0]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[1]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(next_rt_input_router4[2]), .IN2(1'b0), .S(and2result_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U41 ( .A(and2result_input_router4), .Y(invres2_input_router4) );

    AND3X1 U37 ( .IN1(new_rt_input_router4), .IN2(invres1_input_router4), .IN3(invres2_input_router4), .Q(and3result_input_router4) );
    AND2X1 U38 ( .IN1(flit_input_router4[31]), .IN2(1'b1), .Q(and4result_input_router4) );
    AND2X1 U38 ( .IN1(and4result_input_router4), .IN2(and3result_input_router4), .Q(and5result_input_router4) );

    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U38 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[2]);

    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][0]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][1]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][2]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][3]));
    BUFX1 U35(.A(1'sb0), .Y(int_route_v[24:20][4]));

    NOR3X1 U37 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(norres_5_input_router4) );
    AND2X1 U38 ( .IN1(norres_5_input_router4), .IN2(new_rt_input_router4), .Q(and6result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and6result_input_router4), .Q(int_route_v[24:20][4]);

    NOR2X1 U38 ( .IN1(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(and7result_input_router4) );
    AND2X1 U19 ( .IN1(and7result_input_router4), .IN2(next_rt_input_router4[0]), .Y(orres1_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres1_input_router4), .Q(finand1_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router4), .Q(int_route_v[24:20][3]);

    NOR2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[2]), .Q(and8result_input_router4) );
    AND2X1 U19 ( .IN1(and8result_input_router4), .IN2(next_rt_input_router4[1]), .Y(orres2_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres2_input_router4), .Q(finand2_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router4), .Q(int_route_v[24:20][2]);

    NOR2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and9result_input_router4) );
    AND2X1 U19 ( .IN1(and9result_input_router4), .IN2(next_rt_input_router4[2]), .Y(orres3_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(orres3_input_router4), .Q(finand3_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router4), .Q(int_route_v[24:20][0]);

    AND2X1 U38 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and10result_input_router4) );
    INVX1 U41 ( .A(next_rt_input_router4[2]), .Y(nextrt2not_input_router44) );
    AND2X1 U38 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router4), .Q(and11result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    INVX1 U41 ( .A(new_rt_input_router4), .Y(new_rt_input_router4not) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(flit_input_router4_req_i[0]), .Q(secondAndc_input_router4) );

    NOR3X1 U37 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(norres_5_input_router4_2) );
    AND2X1 U38 ( .IN1(norres_5_input_router4_2), .IN2(newsecondAndc_input_router4_rt), .Q(and62result_input_router4) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and62result_input_router4), .Q(int_route_v[24:20][4]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(and7result_input_router42) );
    AND2X1 U19 ( .IN1(and7result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .Y(orres1_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres1_input_router42), .Q(finand1_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router42), .Q(int_route_v[24:20][3]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Q(and8result_input_router42) );
    AND2X1 U19 ( .IN1(and8result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Y(orres2_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres2_input_router4), .Q(finand2_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router42), .Q(int_route_v[24:20][2]);

    NOR2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and9result_input_router42) );
    AND2X1 U19 ( .IN1(and9result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(orres3_input_router42) );
    AND2X1 U38 ( .IN1(new_rt_input_router4not), .IN2(orres3_input_router42), .Q(finand3_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router42), .Q(int_route_v[24:20][0]);

    AND2X1 U38 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and10result_input_router42) );
    INVX1 U41 ( .A(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(nextrt2not_input_router44) );
    AND3X1 U38 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router42), .IN3(new_rt_input_router4not), .Q(and11result_input_router42) );
    MUX21X1 U38 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[0]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[2]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[4]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[5]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[6]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[7]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[8]);
    INVX1 U41 ( .A(arst_value), .Y(arst_valuenot_input_router4) );
    AND2X1 U38 ( .IN1(new_rt_input_router4), .IN2(arst_valuenot_input_router4), .Q(finand3_input_router422) );
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(next_rt_input_router4[0]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(next_rt_input_router4[1]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]);
    MUX21X1 U51 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .IN2(next_rt_input_router4[2]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]); 


//input part


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule[0]), .Y(next_read_ptr_fifomodule[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule[1]), .Y(next_read_ptr_fifomodule[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule[0]), .Y(next_write_ptr_fifomodule[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule[1]), .Y(next_write_ptr_fifomodule[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule[0]), .IN2(read_ptr_ff_fifomodule[0]), .Q(u1temp_fifomodule) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule[1]), .IN2(read_ptr_ff_fifomodule[1]), .Q(u2temp_fifomodule) );
	AND2X1 U3 ( .A(u1temp_fifomodule), .B(u2temp_fifomodule), .Y(empty_vc_buffer) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule[1]), .B(read_ptr_ff_fifomodule[1]), .Y(u4temp_fifomodule) );
	AND2X1 U5 ( .A(u1temp_fifomodule), .B(u4temp_fifomodule), .Y(full_vc_buffer) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][7]));

	INVX1 U7 ( .A(full_vc_buffer), .Y(full_vc_buffer_not_fifomodule) );
	AND2X1 U8 ( .A(write_flit_vc_buffer), .B(full_vc_buffer_not_fifomodule), .Y(u7temp_fifomodule) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule), .Q(u9temp_fifomodule));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule[0]), .B0(u9temp_fifomodule), .C1(u10carry_fifomodule), .SO(next_write_ptr_fifomodule[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule), .B0(write_ptr_ff_fifomodule[1]), .C1(u11carry_fifomodule), .SO(next_write_ptr_fifomodule[1]) );

	INVX1 U12 ( .A(empty_vc_buffer), .Y(empty_vc_buffer_not_fifomodule) );
	AND2X1 U13 ( .A(read_flit_vc_buffer), .B(empty_vc_buffer_not_fifomodule), .Y(u13temp_fifomodule) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule), .Q(u14temp_fifomodule));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule[0]), .B0(u14temp_fifomodule), .C1(u15carry_fifomodule), .SO(next_read_ptr_fifomodule[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule), .B0(read_ptr_ff_fifomodule[1]), .C1(u16carry_fifomodule), .SO(next_read_ptr_fifomodule[1]) );

	AND2X1 U17 ( .A(write_flit_vc_buffer), .B(full_vc_buffer), .Y(u17res_fifomodule) );
	AND2X1 U18 ( .A(read_flit_vc_buffer), .B(empty_vc_buffer), .Y(u18res_fifomodule) );
    OR2X1 U19 ( .A(u17res_fifomodule), .B(u18res_fifomodule), .Y(error_vc_buffer) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule[0]), .B(read_ptr_ff_fifomodule[0]), .Y(fifo_ocup_fifomodule[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule[0]), .Y(write_ptr_ff_fifomodule_0_not) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule_0_not), .B(read_ptr_ff_fifomodule[0]), .Y(b0wire_fifomodule) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule[1]), .B(read_ptr_ff_fifomodule[1]), .Y(u23temp_fifomodule) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule[1]), .Y(write_ptr_ff_fifomodule_1_not) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule[1]), .B(write_ptr_ff_fifomodule_1_not), .Y(boutb_fifomodule) );
	XOR2X1 U24 ( .A(u23temp_fifomodule), .B(b0wire_fifomodule), .Y(fifo_ocup_fifomodule[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule), .Y(u23temp_fifomodule_not_fifomodule) );
	AND2X1 U26 ( .A(b0wire_fifomodule), .B(u23temp_fifomodule_not_fifomodule), .Y(bouta_fifomodule) );
	OR2X1 U27 ( .A(bouta_fifomodule), .B(boutb_fifomodule), .Y(boutmain_fifomodule) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(write_ptr_ff_fifomodule[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(read_ptr_ff_fifomodule[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(fifo_ff_fifomodule[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(write_ptr_ff_fifomodule[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(read_ptr_ff_fifomodule[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(fifo_ff_fifomodule[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule[0]), .Q(write_ptr_ff_fifomodule[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule[1]), .Q(write_ptr_ff_fifomodule[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule[0]), .Q(read_ptr_ff_fifomodule[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule[1]), .Q(read_ptr_ff_fifomodule[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][0]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][1]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][2]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][3]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][4]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][5]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][6]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][7]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer), .Y(next_locked_vc_buffer) );
    BUFX1 U0(.A(flit[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][0]));
	BUFX1 U1(.A(flit[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][1]));
	BUFX1 U2(.A(flit[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][2]));
	BUFX1 U3(.A(flit[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][3]));
	BUFX1 U4(.A(flit[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][4]));
	BUFX1 U5(.A(flit[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][5]));
	BUFX1 U6(.A(flit[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][6]));
	BUFX1 U7(.A(flit[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][7]));
	BUFX1 U8(.A(flit[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][8]));
	BUFX1 U9(.A(flit[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][9]));
	BUFX1 U10(.A(flit[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][10]));
	BUFX1 U11(.A(flit[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][11]));
	BUFX1 U12(.A(flit[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][12]));
	BUFX1 U13(.A(flit[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][13]));
	BUFX1 U14(.A(flit[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][14]));
	BUFX1 U15(.A(flit[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][15]));
	BUFX1 U16(.A(flit[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][16]));
	BUFX1 U17(.A(flit[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][17]));
	BUFX1 U18(.A(flit[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][18]));
	BUFX1 U19(.A(flit[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][19]));
	BUFX1 U20(.A(flit[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][20]));
	BUFX1 U21(.A(flit[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][21]));
	BUFX1 U22(.A(flit[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][22]));
	BUFX1 U23(.A(flit[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][23]));
	BUFX1 U24(.A(flit[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][24]));
	BUFX1 U25(.A(flit[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][25]));
	BUFX1 U26(.A(flit[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][26]));
	BUFX1 U27(.A(flit[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][27]));
	BUFX1 U28(.A(flit[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][28]));
	BUFX1 U29(.A(flit[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][29]));
	BUFX1 U30(.A(flit[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][30]));
	BUFX1 U31(.A(flit[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][31]));
	BUFX1 U32(.A(flit[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][32]));
	BUFX1 U33(.A(flit[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][33]));
    NOR2X1 U34 ( .IN1(flit[33]), .IN2(flit[32]), .QN(norres_vc_buffer_vc_buffer) );
    OR4X1 U35 ( .IN1(flit[29]), .IN2(flit[28]), .IN3(flit[27]), .IN4(flit[26]), .Y(or1res_vc_buffer) );
    OR4X1 U35 ( .IN1(flit[25]), .IN2(flit[24]), .IN3(flit[23]), .IN4(flit[22]), .Y(or2res_vc_buffer) );
    OR2X1 U36 ( .A(or1res_vc_buffer), .B(or2res_vc_buffer), .Y(orres_vc_buffer) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(norres_vc_buffer_vc_buffer), .IN3(orres_vc_buffer), .Q(finres1_vc_buffer) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer), .IN2(1'b1), .S(finres1_vc_buffer), .Q(next_locked_vc_buffer);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(flit[33]), .IN3(flit[32]), .Q(andres1_vc_buffer) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer), .IN2(1'b0), .S(andres1_vc_buffer), .Q(next_locked_vc_buffer);

    INVX1 U41 ( .A(full_vc_buffer), .Y(full_vc_buffer_not) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer), .Y(locked_by_route_ff_vc_buffer_not) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer_not), .S(norres_vc_buffer_vc_buffer), .Q(thirdand_vc_buffer);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(full_vc_buffer_not), .IN3(thirdand_vc_buffer), .Q(write_flit_vc_buffer) );
    AND2X1 U45 ( .IN1(full_vc_buffer_not), .IN2(norres_vc_buffer_vc_buffer), .Q(from_input_resp_input_datapath[0]) );
    INVX1 U46 ( .A(empty_vc_buffer), .Y(to_output_req_in_jump_input_datapathput_datapath[0]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[0]), .IN2(to_output_resp_input_datapath[0]), .Q(read_flit_vc_buffer) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapathput_datapath[2:1]), .Y(2'b00));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer);

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule1[0]), .Y(next_read_ptr_fifomodule1[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule1[1]), .Y(next_read_ptr_fifomodule1[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule1[0]), .Y(next_write_ptr_fifomodule1[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule1[1]), .Y(next_write_ptr_fifomodule1[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule1[0]), .IN2(read_ptr_ff_fifomodule1[0]), .Q(u1temp_fifomodule1) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule1[1]), .IN2(read_ptr_ff_fifomodule1[1]), .Q(u2temp_fifomodule1) );
	AND2X1 U3 ( .A(u1temp_fifomodule1), .B(u2temp_fifomodule1), .Y(empty_vc_buffer1) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule1[1]), .B(read_ptr_ff_fifomodule1[1]), .Y(u4temp_fifomodule1) );
	AND2X1 U5 ( .A(u1temp_fifomodule1), .B(u4temp_fifomodule1), .Y(full_vc_buffer1) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][7]));

	INVX1 U7 ( .A(full_vc_buffer1), .Y(full_vc_buffer1_not1_fifomodule1) );
	AND2X1 U8 ( .A(write_flit1_vc_buffer1), .B(full_vc_buffer1_not1_fifomodule1), .Y(u7temp_fifomodule1) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule1), .Q(u9temp_fifomodule1));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule1[0]), .B0(u9temp_fifomodule1), .C1(u10carry_fifomodule1), .SO(next_write_ptr_fifomodule1[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule1), .B0(write_ptr_ff_fifomodule1[1]), .C1(u11carry_fifomodule1), .SO(next_write_ptr_fifomodule1[1]) );

	INVX1 U12 ( .A(empty_vc_buffer1), .Y(empty_vc_buffer1_not_fifomodule1) );
	AND2X1 U13 ( .A(read_flit1_vc_buffer1), .B(empty_vc_buffer1_not_fifomodule1), .Y(u13temp_fifomodule1) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule1), .Q(u14temp_fifomodule1));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule1[0]), .B0(u14temp_fifomodule1), .C1(u15carry_fifomodule1), .SO(next_read_ptr_fifomodule1[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule1), .B0(read_ptr_ff_fifomodule1[1]), .C1(u16carry_fifomodule1), .SO(next_read_ptr_fifomodule1[1]) );

	AND2X1 U17 ( .A(write_flit1_vc_buffer1), .B(full_vc_buffer1), .Y(u17res_fifomodule1) );
	AND2X1 U18 ( .A(read_flit1_vc_buffer1), .B(empty_vc_buffer1), .Y(u18res_fifomodule1) );
    OR2X1 U19 ( .A(u17res_fifomodule1), .B(u18res_fifomodule1), .Y(error_vc_buffer1) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule1[0]), .B(read_ptr_ff_fifomodule1[0]), .Y(fifo_ocup_fifomodule1[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule1[0]), .Y(write_ptr_ff_fifomodule1_0_not1) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule1_0_not1), .B(read_ptr_ff_fifomodule1[0]), .Y(b0wire_fifomodule1) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule1[1]), .B(read_ptr_ff_fifomodule1[1]), .Y(u23temp_fifomodule1) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule1[1]), .Y(write_ptr_ff_fifomodule1_1_not1) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule1[1]), .B(write_ptr_ff_fifomodule1_1_not1), .Y(boutb_fifomodule1) );
	XOR2X1 U24 ( .A(u23temp_fifomodule1), .B(b0wire_fifomodule1), .Y(fifo_ocup_fifomodule1[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule1), .Y(u23temp_fifomodule1_not_fifomodule1) );
	AND2X1 U26 ( .A(b0wire_fifomodule1), .B(u23temp_fifomodule1_not_fifomodule1), .Y(bouta_fifomodule1) );
	OR2X1 U27 ( .A(bouta_fifomodule1), .B(boutb_fifomodule1), .Y(boutmain_fifomodule1) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule1[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule1[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule1) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule1) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(write_ptr_ff_fifomodule1[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(read_ptr_ff_fifomodule1[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(fifo_ff_fifomodule1[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(write_ptr_ff_fifomodule1[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(read_ptr_ff_fifomodule1[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(fifo_ff_fifomodule1[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule1[0]), .Q(write_ptr_ff_fifomodule1[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule1[1]), .Q(write_ptr_ff_fifomodule1[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule1[0]), .Q(read_ptr_ff_fifomodule1[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule1[1]), .Q(read_ptr_ff_fifomodule1[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][0]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][1]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][2]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][3]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][4]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][5]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][6]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][7]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer1), .Y(next_locked_vc_buffer1) );
    BUFX1 U0(.A(flit1[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][0]));
	BUFX1 U1(.A(flit1[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][1]));
	BUFX1 U2(.A(flit1[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][2]));
	BUFX1 U3(.A(flit1[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][3]));
	BUFX1 U4(.A(flit1[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][4]));
	BUFX1 U5(.A(flit1[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][5]));
	BUFX1 U6(.A(flit1[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][6]));
	BUFX1 U7(.A(flit1[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][7]));
	BUFX1 U8(.A(flit1[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][8]));
	BUFX1 U9(.A(flit1[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][9]));
	BUFX1 U10(.A(flit1[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][10]));
	BUFX1 U11(.A(flit1[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][11]));
	BUFX1 U12(.A(flit1[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][12]));
	BUFX1 U13(.A(flit1[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][13]));
	BUFX1 U14(.A(flit1[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][14]));
	BUFX1 U15(.A(flit1[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][15]));
	BUFX1 U16(.A(flit1[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][16]));
	BUFX1 U17(.A(flit1[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][17]));
	BUFX1 U18(.A(flit1[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][18]));
	BUFX1 U19(.A(flit1[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][19]));
	BUFX1 U20(.A(flit1[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][20]));
	BUFX1 U21(.A(flit1[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][21]));
	BUFX1 U22(.A(flit1[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][22]));
	BUFX1 U23(.A(flit1[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][23]));
	BUFX1 U24(.A(flit1[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][24]));
	BUFX1 U25(.A(flit1[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][25]));
	BUFX1 U26(.A(flit1[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][26]));
	BUFX1 U27(.A(flit1[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][27]));
	BUFX1 U28(.A(flit1[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][28]));
	BUFX1 U29(.A(flit1[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][29]));
	BUFX1 U30(.A(flit1[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][30]));
	BUFX1 U31(.A(flit1[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][31]));
	BUFX1 U32(.A(flit1[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][32]));
	BUFX1 U33(.A(flit1[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][33]));
    NOR2X1 U34 ( .IN1(flit1[33]), .IN2(flit1[32]), .QN(norres_vc_buffer1_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit1[29]), .IN2(flit1[28]), .IN3(flit1[27]), .IN4(flit1[26]), .Y(or1res_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit1[25]), .IN2(flit1[24]), .IN3(flit1[23]), .IN4(flit1[22]), .Y(or2res_vc_buffer1) );
    OR2X1 U36 ( .A(or1res_vc_buffer1), .B(or2res_vc_buffer1), .Y(orres_vc_buffer1) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(norres_vc_buffer1_vc_buffer1), .IN3(orres_vc_buffer1), .Q(finres1_vc_buffer1) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer1), .IN2(1'b1), .S(finres1_vc_buffer1), .Q(next_locked_vc_buffer1);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(flit1[33]), .IN3(flit1[32]), .Q(andres1_vc_buffer1) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer1), .IN2(1'b0), .S(andres1_vc_buffer1), .Q(next_locked_vc_buffer1);

    INVX1 U41 ( .A(full_vc_buffer1), .Y(full_vc_buffer1_not1) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer1), .Y(locked_by_route_ff_vc_buffer1_not1) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer1_not1), .S(norres_vc_buffer1_vc_buffer1), .Q(thirdand_vc_buffer1);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(full_vc_buffer1_not1), .IN3(thirdand_vc_buffer1), .Q(write_flit1_vc_buffer1) );
    AND2X1 U45 ( .IN1(full_vc_buffer1_not1), .IN2(norres_vc_buffer1_vc_buffer1), .Q(from_input_resp_input_datapath[1]) );
    INVX1 U46 ( .A(empty_vc_buffer1), .Y(to_output_req_in_jump_input_datapathput_datapath[37]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[37]), .IN2(to_output_resp_input_datapath[1]), .Q(read_flit1_vc_buffer1) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapathput_datapath[39:38]), .Y(2'b01));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer1), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer1);


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule2[0]), .Y(next_read_ptr_fifomodule2[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule2[1]), .Y(next_read_ptr_fifomodule2[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule2[0]), .Y(next_write_ptr_fifomodule2[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule2[1]), .Y(next_write_ptr_fifomodule2[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule2[0]), .IN2(read_ptr_ff_fifomodule2[0]), .Q(u1temp_fifomodule2) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule2[1]), .IN2(read_ptr_ff_fifomodule2[1]), .Q(u2temp_fifomodule2) );
	AND2X1 U3 ( .A(u1temp_fifomodule2), .B(u2temp_fifomodule2), .Y(empty_vc_buffer2) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule2[1]), .B(read_ptr_ff_fifomodule2[1]), .Y(u4temp_fifomodule2) );
	AND2X1 U5 ( .A(u1temp_fifomodule2), .B(u4temp_fifomodule2), .Y(full_vc_buffer2) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][7]));

	INVX1 U7 ( .A(full_vc_buffer2), .Y(full_vc_buffer2_not2_fifomodule2) );
	AND2X1 U8 ( .A(write_flit2_vc_buffer2), .B(full_vc_buffer2_not2_fifomodule2), .Y(u7temp_fifomodule2) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule2), .Q(u9temp_fifomodule2));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule2[0]), .B0(u9temp_fifomodule2), .C1(u10carry_fifomodule2), .SO(next_write_ptr_fifomodule2[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule2), .B0(write_ptr_ff_fifomodule2[1]), .C1(u11carry_fifomodule2), .SO(next_write_ptr_fifomodule2[1]) );

	INVX1 U12 ( .A(empty_vc_buffer2), .Y(empty_vc_buffer2_not_fifomodule2) );
	AND2X1 U13 ( .A(read_flit2_vc_buffer2), .B(empty_vc_buffer2_not_fifomodule2), .Y(u13temp_fifomodule2) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule2), .Q(u14temp_fifomodule2));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule2[0]), .B0(u14temp_fifomodule2), .C1(u15carry_fifomodule2), .SO(next_read_ptr_fifomodule2[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule2), .B0(read_ptr_ff_fifomodule2[1]), .C1(u16carry_fifomodule2), .SO(next_read_ptr_fifomodule2[1]) );

	AND2X1 U17 ( .A(write_flit2_vc_buffer2), .B(full_vc_buffer2), .Y(u17res_fifomodule2) );
	AND2X1 U18 ( .A(read_flit2_vc_buffer2), .B(empty_vc_buffer2), .Y(u18res_fifomodule2) );
    OR2X1 U19 ( .A(u17res_fifomodule2), .B(u18res_fifomodule2), .Y(error_vc_buffer2) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule2[0]), .B(read_ptr_ff_fifomodule2[0]), .Y(fifo_ocup_fifomodule2[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule2[0]), .Y(write_ptr_ff_fifomodule2_0_not2) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule2_0_not2), .B(read_ptr_ff_fifomodule2[0]), .Y(b0wire_fifomodule2) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule2[1]), .B(read_ptr_ff_fifomodule2[1]), .Y(u23temp_fifomodule2) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule2[1]), .Y(write_ptr_ff_fifomodule2_1_not2) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule2[1]), .B(write_ptr_ff_fifomodule2_1_not2), .Y(boutb_fifomodule2) );
	XOR2X1 U24 ( .A(u23temp_fifomodule2), .B(b0wire_fifomodule2), .Y(fifo_ocup_fifomodule2[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule2), .Y(u23temp_fifomodule2_not_fifomodule2) );
	AND2X1 U26 ( .A(b0wire_fifomodule2), .B(u23temp_fifomodule2_not_fifomodule2), .Y(bouta_fifomodule2) );
	OR2X1 U27 ( .A(bouta_fifomodule2), .B(boutb_fifomodule2), .Y(boutmain_fifomodule2) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule2[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule2[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule2) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule2) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(write_ptr_ff_fifomodule2[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(read_ptr_ff_fifomodule2[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(fifo_ff_fifomodule2[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(write_ptr_ff_fifomodule2[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(read_ptr_ff_fifomodule2[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(fifo_ff_fifomodule2[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule2[0]), .Q(write_ptr_ff_fifomodule2[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule2[1]), .Q(write_ptr_ff_fifomodule2[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule2[0]), .Q(read_ptr_ff_fifomodule2[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule2[1]), .Q(read_ptr_ff_fifomodule2[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][0]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][1]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][2]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][3]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][4]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][5]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][6]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][7]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer2), .Y(next_locked_vc_buffer2) );
    BUFX1 U0(.A(flit2[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][0]));
	BUFX1 U1(.A(flit2[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][1]));
	BUFX1 U2(.A(flit2[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][2]));
	BUFX1 U3(.A(flit2[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][3]));
	BUFX1 U4(.A(flit2[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][4]));
	BUFX1 U5(.A(flit2[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][5]));
	BUFX1 U6(.A(flit2[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][6]));
	BUFX1 U7(.A(flit2[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][7]));
	BUFX1 U8(.A(flit2[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][8]));
	BUFX1 U9(.A(flit2[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][9]));
	BUFX1 U10(.A(flit2[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][10]));
	BUFX1 U11(.A(flit2[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][11]));
	BUFX1 U12(.A(flit2[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][12]));
	BUFX1 U13(.A(flit2[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][13]));
	BUFX1 U14(.A(flit2[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][14]));
	BUFX1 U15(.A(flit2[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][15]));
	BUFX1 U16(.A(flit2[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][16]));
	BUFX1 U17(.A(flit2[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][17]));
	BUFX1 U18(.A(flit2[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][18]));
	BUFX1 U19(.A(flit2[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][19]));
	BUFX1 U20(.A(flit2[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][20]));
	BUFX1 U21(.A(flit2[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][21]));
	BUFX1 U22(.A(flit2[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][22]));
	BUFX1 U23(.A(flit2[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][23]));
	BUFX1 U24(.A(flit2[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][24]));
	BUFX1 U25(.A(flit2[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][25]));
	BUFX1 U26(.A(flit2[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][26]));
	BUFX1 U27(.A(flit2[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][27]));
	BUFX1 U28(.A(flit2[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][28]));
	BUFX1 U29(.A(flit2[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][29]));
	BUFX1 U30(.A(flit2[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][30]));
	BUFX1 U31(.A(flit2[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][31]));
	BUFX1 U32(.A(flit2[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][32]));
	BUFX1 U33(.A(flit2[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][33]));
    NOR2X1 U34 ( .IN1(flit2[33]), .IN2(flit2[32]), .QN(norres_vc_buffer2_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit2[29]), .IN2(flit2[28]), .IN3(flit2[27]), .IN4(flit2[26]), .Y(or1res_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit2[25]), .IN2(flit2[24]), .IN3(flit2[23]), .IN4(flit2[22]), .Y(or2res_vc_buffer2) );
    OR2X1 U36 ( .A(or1res_vc_buffer2), .B(or2res_vc_buffer2), .Y(orres_vc_buffer2) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(norres_vc_buffer2_vc_buffer2), .IN3(orres_vc_buffer2), .Q(finres1_vc_buffer2) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer2), .IN2(1'b1), .S(finres1_vc_buffer2), .Q(next_locked_vc_buffer2);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(flit2[33]), .IN3(flit2[32]), .Q(andres1_vc_buffer2) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer2), .IN2(1'b0), .S(andres1_vc_buffer2), .Q(next_locked_vc_buffer2);

    INVX1 U41 ( .A(full_vc_buffer2), .Y(full_vc_buffer2_not2) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer2), .Y(locked_by_route_ff_vc_buffer2_not2) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer2_not2), .S(norres_vc_buffer2_vc_buffer2), .Q(thirdand_vc_buffer2);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(full_vc_buffer2_not2), .IN3(thirdand_vc_buffer2), .Q(write_flit2_vc_buffer2) );
    AND2X1 U45 ( .IN1(full_vc_buffer2_not2), .IN2(norres_vc_buffer2_vc_buffer2), .Q(from_input_resp_input_datapath[2]) );
    INVX1 U46 ( .A(empty_vc_buffer2), .Y(to_output_req_in_jump_input_datapathput_datapath[74]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[74]), .IN2(to_output_resp_input_datapath[2]), .Q(read_flit2_vc_buffer2) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapathput_datapath[76:75]), .Y(2'b10));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer2), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer2);

	BUFX1 U3(.A(from_input_req_in_jump_input_datapathput_datapath[77]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapathput_datapath[78]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapathput_datapath[79]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapathput_datapath[80]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapathput_datapath[81]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapathput_datapath[82]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapathput_datapath[83]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapathput_datapath[84]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapathput_datapath[85]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapathput_datapath[86]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapathput_datapath[87]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapathput_datapath[88]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapathput_datapath[89]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapathput_datapath[90]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapathput_datapath[91]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapathput_datapath[92]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapathput_datapath[93]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapathput_datapath[94]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapathput_datapath[95]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapathput_datapath[96]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapathput_datapath[97]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapathput_datapath[98]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapathput_datapath[99]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapathput_datapath[100]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapathput_datapath[101]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapathput_datapath[102]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapathput_datapath[103]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapathput_datapath[104]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapathput_datapath[105]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapathput_datapath[106]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapathput_datapath[107]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapathput_datapath[108]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapathput_datapath[109]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapathput_datapath[110]), .Y(ext_req_v_i[36:0][36]));
    XNOR2X1 U222 ( .IN1(ext_req_v_i[36:0][1]), .IN2(i_input_datapath[0]), .QN(xnor1resu_input_datapath) );
    XNOR2X1 U222 ( .IN1(ext_req_v_i[36:0][2]), .IN2(i_input_datapath[1]), .QN(xnor2resu_input_datapath) );
    AND2X1 U128 ( .IN1(xnor1resu_input_datapath), .IN2(xnor2resu_input_datapath), .Q(and1resu_input_datapath) );
    AND3X1 U128 ( .IN1(and1resu_input_datapath), .IN2(ext_req_v_i[36:0][0]), .IN2(ext_req_v_i[36:0][0]), .Q(cond1line_input_datapath) );
    MUX21X1 U0009 (.IN1(vc_ch_act_in_input_datapath[0]), .IN2(i_input_datapath[0]), .S(cond1line_input_datapath), .Q(vc_ch_act_in_input_datapath[0]));
    MUX21X1 U0010 (.IN1(vc_ch_act_in_input_datapath[1]), .IN2(i_input_datapath[1]), .S(cond1line_input_datapath), .Q(vc_ch_act_in_input_datapath[1]));
    MUX21X1 U0011 (.IN1(req_in_jump_input_datapath), .IN2(1), .S(cond1line_input_datapath), .Q(req_in_jump_input_datapath));
	BUFX1 U3(.A(from_input_req_in_jump_input_datapathput_datapath[40]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapathput_datapath[41]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapathput_datapath[42]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapathput_datapath[43]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapathput_datapath[44]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapathput_datapath[45]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapathput_datapath[46]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapathput_datapath[47]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapathput_datapath[48]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapathput_datapath[49]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapathput_datapath[50]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapathput_datapath[51]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapathput_datapath[52]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapathput_datapath[53]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapathput_datapath[54]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapathput_datapath[55]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapathput_datapath[56]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapathput_datapath[57]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapathput_datapath[58]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapathput_datapath[59]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapathput_datapath[60]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapathput_datapath[61]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapathput_datapath[62]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapathput_datapath[63]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapathput_datapath[64]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapathput_datapath[65]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapathput_datapath[66]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapathput_datapath[67]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapathput_datapath[68]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapathput_datapath[69]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapathput_datapath[70]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapathput_datapath[71]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapathput_datapath[72]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapathput_datapath[73]), .Y(ext_req_v_i[36:0][36]));

	BUFX1 U3(.A(from_input_req_in_jump_input_datapathput_datapath[3]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapathput_datapath[4]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapathput_datapath[5]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapathput_datapath[6]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapathput_datapath[7]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapathput_datapath[8]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapathput_datapath[9]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapathput_datapath[10]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapathput_datapath[11]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapathput_datapath[12]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapathput_datapath[13]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapathput_datapath[14]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapathput_datapath[15]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapathput_datapath[16]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapathput_datapath[17]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapathput_datapath[18]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapathput_datapath[19]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapathput_datapath[20]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapathput_datapath[21]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapathput_datapath[22]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapathput_datapath[23]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapathput_datapath[24]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapathput_datapath[25]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapathput_datapath[26]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapathput_datapath[27]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapathput_datapath[28]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapathput_datapath[29]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapathput_datapath[30]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapathput_datapath[31]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapathput_datapath[32]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapathput_datapath[33]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapathput_datapath[34]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapathput_datapath[35]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapathput_datapath[36]), .Y(ext_req_v_i[36:0][36]));

    MUX21X1 U0012 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath * 37]), .IN2(ext_req_v_i[36:0][0]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath * 37]));
    MUX21X1 U0013 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+2]), .IN2(vc_ch_act_in_input_datapath[1]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+2]));
    MUX21X1 U0014 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+1]), .IN2(vc_ch_act_in_input_datapath[0]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+1]));
    MUX21X1 U0015 (.IN1(ext_resp_v_o[1:0][0]), .IN2(from_input_resp_input_datapath[vc_ch_act_in_input_datapath]), .S(req_in_jump_input_datapath), .Q(ext_resp_v_o[1:0][0]));

    INVX1 U041 ( .A(req_in_jump_input_datapath), .Y(req_in_jump_input_datapath_not) );
    MUX21X1 U0016 (.IN1(ext_resp_v_o[1:0][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath_not), .Q(ext_resp_v_o[1:0][0]));
    BUFX1 U34(.A(from_input_req_in_jump_input_datapathput_datapath[34]), .Y(ext_req_v_i[36:0][34]));

    XOR2X1 U0222 ( .IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b1), .Q(xor1resu_input_datapath) );
    MUX21X1 U0017 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(xor1resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U0018 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b0), .S(xor1resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    AND2X1 U38123 ( .IN1(xor1resu_input_datapath), .IN2(to_output_req_in_jump_input_datapathput_datapath[j_input_datapath*37]), .Q(and2resu_input_datapath) );
    MUX21X1 U0019 (.IN1(vc_ch_act_out_input_datapath[0]), .IN2(j_input_datapath[0]), .S(and2resu_input_datapath), .Q(vc_ch_act_out_input_datapath[0]));
    MUX21X1 U0020 (.IN1(vc_ch_act_out_input_datapath[1]), .IN2(j_input_datapath[1]), .S(and2resu_input_datapath), .Q(vc_ch_act_out_input_datapath[1]));
    MUX21X1 U0021 (.IN1(req_out_jump_input_datapath), .IN2(1'b1), .S(and2resu_input_datapath), .Q(req_out_jump_input_datapath));
    MUX21X1 U0022 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(and2resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U0023 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b1), .S(and2resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    HADDX1 U00021 ( .A0(j_input_datapath[0]), .B0(1'b1), .C1(j_input_datapath[1]), .SO(j_input_datapath[0]) );
    HADDX1 U00022 ( .A0(j_input_datapath[0]), .B0(1'b1), .C1(j_input_datapath[1]), .SO(j_input_datapath[0]) );
    AND2X1 U38111 ( .IN1(xor1resu_input_datapath), .IN2(to_output_req_in_jump_input_datapathput_datapath[j_input_datapath*37]), .Q(and3resu) );
    NAND2X1 U29311(.A(_sv2v_jump_input_datapath[0]),.B(_sv2v_jump_input_datapath[1]),.Y(nand1resu_input_datapath));
    MUX21X1 U00212 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(nand1resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U00213 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b0), .S(nand1resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    XNOR2X1 U17581 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(_sv2v_jump_input_datapath[1]), .Q(xnor23resu_input_datapath) );
    AND2X1 U38111 ( .IN1(xnor23resu_input_datapath), .IN2(req_out_jump_input_datapath), .Q(and4resu_input_datapath) );

    MUX21X1 U3(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[36:0][3]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U4(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[36:0][4]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U5(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[36:0][5]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U6(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[36:0][6]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U7(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[36:0][7]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U8(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[36:0][8]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U9(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[36:0][9]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U10(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[36:0][10]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U11(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[36:0][11]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U12(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[36:0][12]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U13(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[36:0][13]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U14(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[36:0][14]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U15(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[36:0][15]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U16(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[36:0][16]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U17(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[36:0][17]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U18(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[36:0][18]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U19(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[36:0][19]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U20(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[36:0][20]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U21(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[36:0][21]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U22(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[36:0][22]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U23(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[36:0][23]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U24(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[36:0][24]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U25(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[36:0][25]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U26(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[36:0][26]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U27(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[36:0][27]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U28(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[36:0][28]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U29(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[36:0][29]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U30(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[36:0][30]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U31(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[36:0][31]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U32(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[36:0][32]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U33(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[36:0][33]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U34(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[36:0][34]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U35(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[36:0][35]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U36(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[36:0][36]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U321111(.IN1(int_req_v[36:0][0]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath * 37)]), .S(and4resu_input_datapath), .Q(int_req_v[36:0][0]));
	MUX21X1 U331112(.IN1(int_req_v[36:0][1]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+1]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+1]));
	MUX21X1 U331122(.IN1(int_req_v[36:0][2]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+2]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath[vc_ch_act_out_input_datapath]),.IN2(int_resp_v[1:0]), .S(and4resu_input_datapath), .Q(to_output_resp_input_datapath[vc_ch_act_out_input_datapath]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath[vc_ch_act_out_input_datapath+1]),.IN2(int_resp_v[1:0]), .S(and4resu_input_datapath), .Q(to_output_resp_input_datapath[vc_ch_act_out_input_datapath+1]));


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule11[0]), .Y(next_read_ptr_fifomodule11[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule11[1]), .Y(next_read_ptr_fifomodule11[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule11[0]), .Y(next_write_ptr_fifomodule11[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule11[1]), .Y(next_write_ptr_fifomodule11[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule11[0]), .IN2(read_ptr_ff_fifomodule11[0]), .Q(u1temp_fifomodule11) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule11[1]), .IN2(read_ptr_ff_fifomodule11[1]), .Q(u2temp_fifomodule11) );
	AND2X1 U3 ( .A(u1temp_fifomodule11), .B(u2temp_fifomodule11), .Y(empty_vc_buffer11) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule11[1]), .B(read_ptr_ff_fifomodule11[1]), .Y(u4temp_fifomodule11) );
	AND2X1 U5 ( .A(u1temp_fifomodule11), .B(u4temp_fifomodule11), .Y(full_vc_buffer11) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][7]));

	INVX1 U7 ( .A(full_vc_buffer11), .Y(full_vc_buffer11_not_fifomodule) );
	AND2X1 U8 ( .A(write_flit11_vc_buffer1), .B(full_vc_buffer11_not_fifomodule), .Y(u7temp_fifomodule11) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule11), .Q(u9temp_fifomodule11));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule11[0]), .B0(u9temp_fifomodule11), .C1(u10carry_fifomodule11), .SO(next_write_ptr_fifomodule11[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule11), .B0(write_ptr_ff_fifomodule11[1]), .C1(u11carry_fifomodule11), .SO(next_write_ptr_fifomodule11[1]) );

	INVX1 U12 ( .A(empty_vc_buffer11), .Y(empty_vc_buffer11_not_fifomodule) );
	AND2X1 U13 ( .A(read_flit11_vc_buffer1), .B(empty_vc_buffer11_not_fifomodule), .Y(u13temp_fifomodule11) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule11), .Q(u14temp_fifomodule11));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule11[0]), .B0(u14temp_fifomodule11), .C1(u15carry_fifomodule11), .SO(next_read_ptr_fifomodule11[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule11), .B0(read_ptr_ff_fifomodule11[1]), .C1(u16carry_fifomodule11), .SO(next_read_ptr_fifomodule11[1]) );

	AND2X1 U17 ( .A(write_flit11_vc_buffer1), .B(full_vc_buffer11), .Y(u17res_fifomodule11) );
	AND2X1 U18 ( .A(read_flit11_vc_buffer1), .B(empty_vc_buffer11), .Y(u18res_fifomodule11) );
    OR2X1 U19 ( .A(u17res_fifomodule11), .B(u18res_fifomodule11), .Y(error_vc_buffer11) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule11[0]), .B(read_ptr_ff_fifomodule11[0]), .Y(fifo_ocup_fifomodule11[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule11[0]), .Y(write_ptr_ff_fifomodule11_0_not1) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule11_0_not1), .B(read_ptr_ff_fifomodule11[0]), .Y(b0wire_fifomodule11) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule11[1]), .B(read_ptr_ff_fifomodule11[1]), .Y(u23temp_fifomodule11) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule11[1]), .Y(write_ptr_ff_fifomodule11_1_not1) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule11[1]), .B(write_ptr_ff_fifomodule11_1_not1), .Y(boutb_fifomodule11) );
	XOR2X1 U24 ( .A(u23temp_fifomodule11), .B(b0wire_fifomodule11), .Y(fifo_ocup_fifomodule11[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule11), .Y(u23temp_fifomodule11_not_fifomodule11) );
	AND2X1 U26 ( .A(b0wire_fifomodule11), .B(u23temp_fifomodule11_not_fifomodule11), .Y(bouta_fifomodule11) );
	OR2X1 U27 ( .A(bouta_fifomodule11), .B(boutb_fifomodule11), .Y(boutmain_fifomodule11) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule11[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule11[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule11) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule11) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(write_ptr_ff_fifomodule11[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(read_ptr_ff_fifomodule11[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(fifo_ff_fifomodule11[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(write_ptr_ff_fifomodule11[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(read_ptr_ff_fifomodule11[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(fifo_ff_fifomodule11[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule11[0]), .Q(write_ptr_ff_fifomodule11[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule11[1]), .Q(write_ptr_ff_fifomodule11[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule11[0]), .Q(read_ptr_ff_fifomodule11[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule11[1]), .Q(read_ptr_ff_fifomodule11[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][0]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][1]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][2]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][3]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][4]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][5]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][6]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][7]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer11), .Y(next_locked_vc_buffer11) );
    BUFX1 U0(.A(flit11[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][0]));
	BUFX1 U1(.A(flit11[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][1]));
	BUFX1 U2(.A(flit11[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][2]));
	BUFX1 U3(.A(flit11[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][3]));
	BUFX1 U4(.A(flit11[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][4]));
	BUFX1 U5(.A(flit11[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][5]));
	BUFX1 U6(.A(flit11[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][6]));
	BUFX1 U7(.A(flit11[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][7]));
	BUFX1 U8(.A(flit11[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][8]));
	BUFX1 U9(.A(flit11[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][9]));
	BUFX1 U10(.A(flit11[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][10]));
	BUFX1 U11(.A(flit11[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][11]));
	BUFX1 U12(.A(flit11[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][12]));
	BUFX1 U13(.A(flit11[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][13]));
	BUFX1 U14(.A(flit11[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][14]));
	BUFX1 U15(.A(flit11[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][15]));
	BUFX1 U16(.A(flit11[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][16]));
	BUFX1 U17(.A(flit11[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][17]));
	BUFX1 U18(.A(flit11[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][18]));
	BUFX1 U19(.A(flit11[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][19]));
	BUFX1 U20(.A(flit11[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][20]));
	BUFX1 U21(.A(flit11[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][21]));
	BUFX1 U22(.A(flit11[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][22]));
	BUFX1 U23(.A(flit11[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][23]));
	BUFX1 U24(.A(flit11[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][24]));
	BUFX1 U25(.A(flit11[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][25]));
	BUFX1 U26(.A(flit11[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][26]));
	BUFX1 U27(.A(flit11[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][27]));
	BUFX1 U28(.A(flit11[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][28]));
	BUFX1 U29(.A(flit11[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][29]));
	BUFX1 U30(.A(flit11[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][30]));
	BUFX1 U31(.A(flit11[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][31]));
	BUFX1 U32(.A(flit11[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][32]));
	BUFX1 U33(.A(flit11[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][33]));
    NOR2X1 U34 ( .IN1(flit11[33]), .IN2(flit11[32]), .QN(norres_vc_buffer11_vc_buffer11) );
    OR4X1 U35 ( .IN1(flit11[29]), .IN2(flit11[28]), .IN3(flit11[27]), .IN4(flit11[26]), .Y(or1res_vc_buffer11) );
    OR4X1 U35 ( .IN1(flit11[25]), .IN2(flit11[24]), .IN3(flit11[23]), .IN4(flit11[22]), .Y(or2res_vc_buffer11) );
    OR2X1 U36 ( .A(or1res_vc_buffer11), .B(or2res_vc_buffer11), .Y(orres_vc_buffer11) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(norres_vc_buffer11_vc_buffer11), .IN3(orres_vc_buffer11), .Q(finres1_vc_buffer11) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer11), .IN2(1'b1), .S(finres1_vc_buffer11), .Q(next_locked_vc_buffer11);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(flit11[33]), .IN3(flit11[32]), .Q(andres1_vc_buffer11) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer11), .IN2(1'b0), .S(andres1_vc_buffer11), .Q(next_locked_vc_buffer11);

    INVX1 U41 ( .A(full_vc_buffer11), .Y(full_vc_buffer11_not) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer11), .Y(locked_by_route_ff_vc_buffer11_not) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer11_not), .S(norres_vc_buffer11_vc_buffer11), .Q(thirdand_vc_buffer11);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(full_vc_buffer11_not), .IN3(thirdand_vc_buffer11), .Q(write_flit11_vc_buffer1) );
    AND2X1 U45 ( .IN1(full_vc_buffer11_not), .IN2(norres_vc_buffer11_vc_buffer11), .Q(from_input_resp_input_datapath1[0]) );
    INVX1 U46 ( .A(empty_vc_buffer11), .Y(to_output_req_in_jump_input_datapath1put_datapath1[0]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[0]), .IN2(to_output_resp_input_datapath1[0]), .Q(read_flit11_vc_buffer1) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath1put_datapath1[2:1]), .Y(2'b00));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer11), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer11);

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule111[0]), .Y(next_read_ptr_fifomodule111[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule111[1]), .Y(next_read_ptr_fifomodule111[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule111[0]), .Y(next_write_ptr_fifomodule111[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule111[1]), .Y(next_write_ptr_fifomodule111[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule111[0]), .IN2(read_ptr_ff_fifomodule111[0]), .Q(u1temp_fifomodule111) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule111[1]), .IN2(read_ptr_ff_fifomodule111[1]), .Q(u2temp_fifomodule111) );
	AND2X1 U3 ( .A(u1temp_fifomodule111), .B(u2temp_fifomodule111), .Y(empty_vc_buffer111) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule111[1]), .B(read_ptr_ff_fifomodule111[1]), .Y(u4temp_fifomodule111) );
	AND2X1 U5 ( .A(u1temp_fifomodule111), .B(u4temp_fifomodule111), .Y(full_vc_buffer111) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][7]));

	INVX1 U7 ( .A(full_vc_buffer111), .Y(full_vc_buffer111_not1_fifomodule1) );
	AND2X1 U8 ( .A(write_flit111_vc_buffer11), .B(full_vc_buffer111_not1_fifomodule1), .Y(u7temp_fifomodule111) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule111), .Q(u9temp_fifomodule111));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule111[0]), .B0(u9temp_fifomodule111), .C1(u10carry_fifomodule111), .SO(next_write_ptr_fifomodule111[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule111), .B0(write_ptr_ff_fifomodule111[1]), .C1(u11carry_fifomodule111), .SO(next_write_ptr_fifomodule111[1]) );

	INVX1 U12 ( .A(empty_vc_buffer111), .Y(empty_vc_buffer111_not_fifomodule1) );
	AND2X1 U13 ( .A(read_flit111_vc_buffer11), .B(empty_vc_buffer111_not_fifomodule1), .Y(u13temp_fifomodule111) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule111), .Q(u14temp_fifomodule111));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule111[0]), .B0(u14temp_fifomodule111), .C1(u15carry_fifomodule111), .SO(next_read_ptr_fifomodule111[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule111), .B0(read_ptr_ff_fifomodule111[1]), .C1(u16carry_fifomodule111), .SO(next_read_ptr_fifomodule111[1]) );

	AND2X1 U17 ( .A(write_flit111_vc_buffer11), .B(full_vc_buffer111), .Y(u17res_fifomodule111) );
	AND2X1 U18 ( .A(read_flit111_vc_buffer11), .B(empty_vc_buffer111), .Y(u18res_fifomodule111) );
    OR2X1 U19 ( .A(u17res_fifomodule111), .B(u18res_fifomodule111), .Y(error_vc_buffer111) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule111[0]), .B(read_ptr_ff_fifomodule111[0]), .Y(fifo_ocup_fifomodule111[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule111[0]), .Y(write_ptr_ff_fifomodule111_0_not11) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule111_0_not11), .B(read_ptr_ff_fifomodule111[0]), .Y(b0wire_fifomodule111) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule111[1]), .B(read_ptr_ff_fifomodule111[1]), .Y(u23temp_fifomodule111) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule111[1]), .Y(write_ptr_ff_fifomodule111_1_not11) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule111[1]), .B(write_ptr_ff_fifomodule111_1_not11), .Y(boutb_fifomodule111) );
	XOR2X1 U24 ( .A(u23temp_fifomodule111), .B(b0wire_fifomodule111), .Y(fifo_ocup_fifomodule111[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule111), .Y(u23temp_fifomodule111_not_fifomodule1) );
	AND2X1 U26 ( .A(b0wire_fifomodule111), .B(u23temp_fifomodule111_not_fifomodule1), .Y(bouta_fifomodule111) );
	OR2X1 U27 ( .A(bouta_fifomodule111), .B(boutb_fifomodule111), .Y(boutmain_fifomodule111) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule111[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule111[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule111) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule111) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(write_ptr_ff_fifomodule111[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(read_ptr_ff_fifomodule111[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(fifo_ff_fifomodule111[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(write_ptr_ff_fifomodule111[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(read_ptr_ff_fifomodule111[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(fifo_ff_fifomodule111[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule111[0]), .Q(write_ptr_ff_fifomodule111[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule111[1]), .Q(write_ptr_ff_fifomodule111[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule111[0]), .Q(read_ptr_ff_fifomodule111[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule111[1]), .Q(read_ptr_ff_fifomodule111[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][0]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][1]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][2]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][3]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][4]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][5]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][6]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][7]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer111), .Y(next_locked_vc_buffer111) );
    BUFX1 U0(.A(flit111[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][0]));
	BUFX1 U1(.A(flit111[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][1]));
	BUFX1 U2(.A(flit111[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][2]));
	BUFX1 U3(.A(flit111[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][3]));
	BUFX1 U4(.A(flit111[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][4]));
	BUFX1 U5(.A(flit111[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][5]));
	BUFX1 U6(.A(flit111[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][6]));
	BUFX1 U7(.A(flit111[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][7]));
	BUFX1 U8(.A(flit111[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][8]));
	BUFX1 U9(.A(flit111[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][9]));
	BUFX1 U10(.A(flit111[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][10]));
	BUFX1 U11(.A(flit111[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][11]));
	BUFX1 U12(.A(flit111[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][12]));
	BUFX1 U13(.A(flit111[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][13]));
	BUFX1 U14(.A(flit111[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][14]));
	BUFX1 U15(.A(flit111[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][15]));
	BUFX1 U16(.A(flit111[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][16]));
	BUFX1 U17(.A(flit111[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][17]));
	BUFX1 U18(.A(flit111[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][18]));
	BUFX1 U19(.A(flit111[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][19]));
	BUFX1 U20(.A(flit111[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][20]));
	BUFX1 U21(.A(flit111[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][21]));
	BUFX1 U22(.A(flit111[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][22]));
	BUFX1 U23(.A(flit111[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][23]));
	BUFX1 U24(.A(flit111[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][24]));
	BUFX1 U25(.A(flit111[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][25]));
	BUFX1 U26(.A(flit111[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][26]));
	BUFX1 U27(.A(flit111[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][27]));
	BUFX1 U28(.A(flit111[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][28]));
	BUFX1 U29(.A(flit111[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][29]));
	BUFX1 U30(.A(flit111[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][30]));
	BUFX1 U31(.A(flit111[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][31]));
	BUFX1 U32(.A(flit111[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][32]));
	BUFX1 U33(.A(flit111[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][33]));
    NOR2X1 U34 ( .IN1(flit111[33]), .IN2(flit111[32]), .QN(norres_vc_buffer111_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit111[29]), .IN2(flit111[28]), .IN3(flit111[27]), .IN4(flit111[26]), .Y(or1res_vc_buffer111) );
    OR4X1 U35 ( .IN1(flit111[25]), .IN2(flit111[24]), .IN3(flit111[23]), .IN4(flit111[22]), .Y(or2res_vc_buffer111) );
    OR2X1 U36 ( .A(or1res_vc_buffer111), .B(or2res_vc_buffer111), .Y(orres_vc_buffer111) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(norres_vc_buffer111_vc_buffer1), .IN3(orres_vc_buffer111), .Q(finres1_vc_buffer111) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer111), .IN2(1'b1), .S(finres1_vc_buffer111), .Q(next_locked_vc_buffer111);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(flit111[33]), .IN3(flit111[32]), .Q(andres1_vc_buffer111) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer111), .IN2(1'b0), .S(andres1_vc_buffer111), .Q(next_locked_vc_buffer111);

    INVX1 U41 ( .A(full_vc_buffer111), .Y(full_vc_buffer111_not1) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer111), .Y(locked_by_route_ff_vc_buffer111_not1) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer111_not1), .S(norres_vc_buffer111_vc_buffer1), .Q(thirdand_vc_buffer111);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(full_vc_buffer111_not1), .IN3(thirdand_vc_buffer111), .Q(write_flit111_vc_buffer11) );
    AND2X1 U45 ( .IN1(full_vc_buffer111_not1), .IN2(norres_vc_buffer111_vc_buffer1), .Q(from_input_resp_input_datapath1[1]) );
    INVX1 U46 ( .A(empty_vc_buffer111), .Y(to_output_req_in_jump_input_datapath1put_datapath1[37]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[37]), .IN2(to_output_resp_input_datapath1[1]), .Q(read_flit111_vc_buffer11) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath1put_datapath1[39:38]), .Y(2'b01));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer111), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer111);


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule112[0]), .Y(next_read_ptr_fifomodule112[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule112[1]), .Y(next_read_ptr_fifomodule112[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule112[0]), .Y(next_write_ptr_fifomodule112[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule112[1]), .Y(next_write_ptr_fifomodule112[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule112[0]), .IN2(read_ptr_ff_fifomodule112[0]), .Q(u1temp_fifomodule112) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule112[1]), .IN2(read_ptr_ff_fifomodule112[1]), .Q(u2temp_fifomodule112) );
	AND2X1 U3 ( .A(u1temp_fifomodule112), .B(u2temp_fifomodule112), .Y(empty_vc_buffer112) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule112[1]), .B(read_ptr_ff_fifomodule112[1]), .Y(u4temp_fifomodule112) );
	AND2X1 U5 ( .A(u1temp_fifomodule112), .B(u4temp_fifomodule112), .Y(full_vc_buffer112) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][7]));

	INVX1 U7 ( .A(full_vc_buffer112), .Y(full_vc_buffer112_not2_fifomodule2) );
	AND2X1 U8 ( .A(write_flit112_vc_buffer21), .B(full_vc_buffer112_not2_fifomodule2), .Y(u7temp_fifomodule112) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule112), .Q(u9temp_fifomodule112));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule112[0]), .B0(u9temp_fifomodule112), .C1(u10carry_fifomodule112), .SO(next_write_ptr_fifomodule112[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule112), .B0(write_ptr_ff_fifomodule112[1]), .C1(u11carry_fifomodule112), .SO(next_write_ptr_fifomodule112[1]) );

	INVX1 U12 ( .A(empty_vc_buffer112), .Y(empty_vc_buffer112_not_fifomodule2) );
	AND2X1 U13 ( .A(read_flit112_vc_buffer21), .B(empty_vc_buffer112_not_fifomodule2), .Y(u13temp_fifomodule112) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule112), .Q(u14temp_fifomodule112));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule112[0]), .B0(u14temp_fifomodule112), .C1(u15carry_fifomodule112), .SO(next_read_ptr_fifomodule112[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule112), .B0(read_ptr_ff_fifomodule112[1]), .C1(u16carry_fifomodule112), .SO(next_read_ptr_fifomodule112[1]) );

	AND2X1 U17 ( .A(write_flit112_vc_buffer21), .B(full_vc_buffer112), .Y(u17res_fifomodule112) );
	AND2X1 U18 ( .A(read_flit112_vc_buffer21), .B(empty_vc_buffer112), .Y(u18res_fifomodule112) );
    OR2X1 U19 ( .A(u17res_fifomodule112), .B(u18res_fifomodule112), .Y(error_vc_buffer112) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule112[0]), .B(read_ptr_ff_fifomodule112[0]), .Y(fifo_ocup_fifomodule112[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule112[0]), .Y(write_ptr_ff_fifomodule112_0_not21) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule112_0_not21), .B(read_ptr_ff_fifomodule112[0]), .Y(b0wire_fifomodule112) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule112[1]), .B(read_ptr_ff_fifomodule112[1]), .Y(u23temp_fifomodule112) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule112[1]), .Y(write_ptr_ff_fifomodule112_1_not21) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule112[1]), .B(write_ptr_ff_fifomodule112_1_not21), .Y(boutb_fifomodule112) );
	XOR2X1 U24 ( .A(u23temp_fifomodule112), .B(b0wire_fifomodule112), .Y(fifo_ocup_fifomodule112[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule112), .Y(u23temp_fifomodule112_not_fifomodule2) );
	AND2X1 U26 ( .A(b0wire_fifomodule112), .B(u23temp_fifomodule112_not_fifomodule2), .Y(bouta_fifomodule112) );
	OR2X1 U27 ( .A(bouta_fifomodule112), .B(boutb_fifomodule112), .Y(boutmain_fifomodule112) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule112[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule112[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule112) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule112) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(write_ptr_ff_fifomodule112[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(read_ptr_ff_fifomodule112[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(fifo_ff_fifomodule112[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(write_ptr_ff_fifomodule112[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(read_ptr_ff_fifomodule112[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(fifo_ff_fifomodule112[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule112[0]), .Q(write_ptr_ff_fifomodule112[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule112[1]), .Q(write_ptr_ff_fifomodule112[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule112[0]), .Q(read_ptr_ff_fifomodule112[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule112[1]), .Q(read_ptr_ff_fifomodule112[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][0]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][1]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][2]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][3]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][4]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][5]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][6]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][7]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer112), .Y(next_locked_vc_buffer112) );
    BUFX1 U0(.A(flit112[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][0]));
	BUFX1 U1(.A(flit112[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][1]));
	BUFX1 U2(.A(flit112[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][2]));
	BUFX1 U3(.A(flit112[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][3]));
	BUFX1 U4(.A(flit112[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][4]));
	BUFX1 U5(.A(flit112[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][5]));
	BUFX1 U6(.A(flit112[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][6]));
	BUFX1 U7(.A(flit112[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][7]));
	BUFX1 U8(.A(flit112[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][8]));
	BUFX1 U9(.A(flit112[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][9]));
	BUFX1 U10(.A(flit112[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][10]));
	BUFX1 U11(.A(flit112[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][11]));
	BUFX1 U12(.A(flit112[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][12]));
	BUFX1 U13(.A(flit112[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][13]));
	BUFX1 U14(.A(flit112[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][14]));
	BUFX1 U15(.A(flit112[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][15]));
	BUFX1 U16(.A(flit112[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][16]));
	BUFX1 U17(.A(flit112[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][17]));
	BUFX1 U18(.A(flit112[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][18]));
	BUFX1 U19(.A(flit112[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][19]));
	BUFX1 U20(.A(flit112[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][20]));
	BUFX1 U21(.A(flit112[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][21]));
	BUFX1 U22(.A(flit112[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][22]));
	BUFX1 U23(.A(flit112[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][23]));
	BUFX1 U24(.A(flit112[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][24]));
	BUFX1 U25(.A(flit112[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][25]));
	BUFX1 U26(.A(flit112[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][26]));
	BUFX1 U27(.A(flit112[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][27]));
	BUFX1 U28(.A(flit112[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][28]));
	BUFX1 U29(.A(flit112[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][29]));
	BUFX1 U30(.A(flit112[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][30]));
	BUFX1 U31(.A(flit112[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][31]));
	BUFX1 U32(.A(flit112[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][32]));
	BUFX1 U33(.A(flit112[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][33]));
    NOR2X1 U34 ( .IN1(flit112[33]), .IN2(flit112[32]), .QN(norres_vc_buffer112_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit112[29]), .IN2(flit112[28]), .IN3(flit112[27]), .IN4(flit112[26]), .Y(or1res_vc_buffer112) );
    OR4X1 U35 ( .IN1(flit112[25]), .IN2(flit112[24]), .IN3(flit112[23]), .IN4(flit112[22]), .Y(or2res_vc_buffer112) );
    OR2X1 U36 ( .A(or1res_vc_buffer112), .B(or2res_vc_buffer112), .Y(orres_vc_buffer112) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(norres_vc_buffer112_vc_buffer2), .IN3(orres_vc_buffer112), .Q(finres1_vc_buffer112) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer112), .IN2(1'b1), .S(finres1_vc_buffer112), .Q(next_locked_vc_buffer112);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(flit112[33]), .IN3(flit112[32]), .Q(andres1_vc_buffer112) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer112), .IN2(1'b0), .S(andres1_vc_buffer112), .Q(next_locked_vc_buffer112);

    INVX1 U41 ( .A(full_vc_buffer112), .Y(full_vc_buffer112_not2) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer112), .Y(locked_by_route_ff_vc_buffer112_not2) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer112_not2), .S(norres_vc_buffer112_vc_buffer2), .Q(thirdand_vc_buffer112);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(full_vc_buffer112_not2), .IN3(thirdand_vc_buffer112), .Q(write_flit112_vc_buffer21) );
    AND2X1 U45 ( .IN1(full_vc_buffer112_not2), .IN2(norres_vc_buffer112_vc_buffer2), .Q(from_input_resp_input_datapath1[2]) );
    INVX1 U46 ( .A(empty_vc_buffer112), .Y(to_output_req_in_jump_input_datapath1put_datapath1[74]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[74]), .IN2(to_output_resp_input_datapath1[2]), .Q(read_flit112_vc_buffer21) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath1put_datapath1[76:75]), .Y(2'b10));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer112), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer112);

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath1put_datapath1[77]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath1put_datapath1[78]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath1put_datapath1[79]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath1put_datapath1[80]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath1put_datapath1[81]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath1put_datapath1[82]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath1put_datapath1[83]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath1put_datapath1[84]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath1put_datapath1[85]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath1put_datapath1[86]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath1put_datapath1[87]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath1put_datapath1[88]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath1put_datapath1[89]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath1put_datapath1[90]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath1put_datapath1[91]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath1put_datapath1[92]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath1put_datapath1[93]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath1put_datapath1[94]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath1put_datapath1[95]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath1put_datapath1[96]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath1put_datapath1[97]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath1put_datapath1[98]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath1put_datapath1[99]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath1put_datapath1[100]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath1put_datapath1[101]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath1put_datapath1[102]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath1put_datapath1[103]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath1put_datapath1[104]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath1put_datapath1[105]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath1put_datapath1[106]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath1put_datapath1[107]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath1put_datapath1[108]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath1put_datapath1[109]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath1put_datapath1[110]), .Y(ext_req_v_i[73:37][36]));
    XNOR2X1 U222 ( .IN1(ext_req_v_i[73:37][1]), .IN2(i_input_datapath1[0]), .QN(xnor1resu_input_datapath1) );
    XNOR2X1 U222 ( .IN1(ext_req_v_i[73:37][2]), .IN2(i_input_datapath1[1]), .QN(xnor2resu_input_datapath1) );
    AND2X1 U128 ( .IN1(xnor1resu_input_datapath1), .IN2(xnor2resu_input_datapath1), .Q(and1resu_input_datapath1) );
    AND3X1 U128 ( .IN1(and1resu_input_datapath1), .IN2(ext_req_v_i[73:37][0]), .IN2(ext_req_v_i[73:37][0]), .Q(cond1line_input_datapath1) );
    MUX21X1 U0009 (.IN1(vc_ch_act_in_input_datapath1[0]), .IN2(i_input_datapath1[0]), .S(cond1line_input_datapath1), .Q(vc_ch_act_in_input_datapath1[0]));
    MUX21X1 U0010 (.IN1(vc_ch_act_in_input_datapath1[1]), .IN2(i_input_datapath1[1]), .S(cond1line_input_datapath1), .Q(vc_ch_act_in_input_datapath1[1]));
    MUX21X1 U0011 (.IN1(req_in_jump_input_datapath1), .IN2(1), .S(cond1line_input_datapath1), .Q(req_in_jump_input_datapath1));
	BUFX1 U3(.A(from_input_req_in_jump_input_datapath1put_datapath1[40]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath1put_datapath1[41]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath1put_datapath1[42]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath1put_datapath1[43]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath1put_datapath1[44]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath1put_datapath1[45]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath1put_datapath1[46]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath1put_datapath1[47]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath1put_datapath1[48]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath1put_datapath1[49]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath1put_datapath1[50]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath1put_datapath1[51]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath1put_datapath1[52]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath1put_datapath1[53]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath1put_datapath1[54]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath1put_datapath1[55]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath1put_datapath1[56]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath1put_datapath1[57]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath1put_datapath1[58]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath1put_datapath1[59]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath1put_datapath1[60]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath1put_datapath1[61]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath1put_datapath1[62]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath1put_datapath1[63]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath1put_datapath1[64]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath1put_datapath1[65]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath1put_datapath1[66]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath1put_datapath1[67]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath1put_datapath1[68]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath1put_datapath1[69]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath1put_datapath1[70]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath1put_datapath1[71]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath1put_datapath1[72]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath1put_datapath1[73]), .Y(ext_req_v_i[73:37][36]));

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath1put_datapath1[3]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath1put_datapath1[4]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath1put_datapath1[5]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath1put_datapath1[6]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath1put_datapath1[7]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath1put_datapath1[8]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath1put_datapath1[9]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath1put_datapath1[10]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath1put_datapath1[11]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath1put_datapath1[12]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath1put_datapath1[13]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath1put_datapath1[14]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath1put_datapath1[15]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath1put_datapath1[16]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath1put_datapath1[17]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath1put_datapath1[18]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath1put_datapath1[19]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath1put_datapath1[20]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath1put_datapath1[21]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath1put_datapath1[22]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath1put_datapath1[23]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath1put_datapath1[24]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath1put_datapath1[25]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath1put_datapath1[26]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath1put_datapath1[27]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath1put_datapath1[28]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath1put_datapath1[29]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath1put_datapath1[30]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath1put_datapath1[31]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath1put_datapath1[32]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath1put_datapath1[33]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath1put_datapath1[34]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath1put_datapath1[35]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath1put_datapath1[36]), .Y(ext_req_v_i[73:37][36]));

    MUX21X1 U0012 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1 * 37]), .IN2(ext_req_v_i[73:37][0]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1 * 37]));
    MUX21X1 U0013 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+2]), .IN2(vc_ch_act_in_input_datapath1[1]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+2]));
    MUX21X1 U0014 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+1]), .IN2(vc_ch_act_in_input_datapath1[0]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+1]));
    MUX21X1 U0015 (.IN1(ext_resp_v_o[2:1][0]), .IN2(from_input_resp_input_datapath1[vc_ch_act_in_input_datapath1]), .S(req_in_jump_input_datapath1), .Q(ext_resp_v_o[2:1][0]));

    INVX1 U041 ( .A(req_in_jump_input_datapath1), .Y(req_in_jump_input_datapath1_not) );
    MUX21X1 U0016 (.IN1(ext_resp_v_o[2:1][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath1_not), .Q(ext_resp_v_o[2:1][0]));
    BUFX1 U34(.A(from_input_req_in_jump_input_datapath1put_datapath1[34]), .Y(ext_req_v_i[73:37][34]));

    XOR2X1 U0222 ( .IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b1), .Q(xor1resu_input_datapath1) );
    MUX21X1 U0017 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(xor1resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U0018 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b0), .S(xor1resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[1]));
    AND2X1 U38123 ( .IN1(xor1resu_input_datapath1), .IN2(to_output_req_in_jump_input_datapath1put_datapath1[j_input_datapath1*37]), .Q(and2resu_input_datapath1) );
    MUX21X1 U0019 (.IN1(vc_ch_act_out_input_datapath1[0]), .IN2(j_input_datapath1[0]), .S(and2resu_input_datapath1), .Q(vc_ch_act_out_input_datapath1[0]));
    MUX21X1 U0020 (.IN1(vc_ch_act_out_input_datapath1[1]), .IN2(j_input_datapath1[1]), .S(and2resu_input_datapath1), .Q(vc_ch_act_out_input_datapath1[1]));
    MUX21X1 U0021 (.IN1(req_out_jump_input_datapath1), .IN2(1'b1), .S(and2resu_input_datapath1), .Q(req_out_jump_input_datapath1));
    MUX21X1 U0022 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(and2resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U0023 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b1), .S(and2resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[1]));
    HADDX1 U00021 ( .A0(j_input_datapath1[0]), .B0(1'b1), .C1(j_input_datapath1[1]), .SO(j_input_datapath1[0]) );
    HADDX1 U00022 ( .A0(j_input_datapath1[0]), .B0(1'b1), .C1(j_input_datapath1[1]), .SO(j_input_datapath1[0]) );
    AND2X1 U38111 ( .IN1(xor1resu_input_datapath1), .IN2(to_output_req_in_jump_input_datapath1put_datapath1[j_input_datapath1*37]), .Q(and3resu) );
    NAND2X1 U29311(.A(_sv2v_jump_input_datapath1[0]),.B(_sv2v_jump_input_datapath1[1]),.Y(nand1resu_input_datapath11));
    MUX21X1 U00212 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(nand1resu_input_datapath11), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U00213 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b0), .S(nand1resu_input_datapath11), .Q(_sv2v_jump_input_datapath1[1]));
    XNOR2X1 U17581 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(_sv2v_jump_input_datapath1[1]), .Q(xnor23resu_input_datapath1) );
    AND2X1 U38111 ( .IN1(xnor23resu_input_datapath1), .IN2(req_out_jump_input_datapath1), .Q(and4resu_input_datapath1) );

    MUX21X1 U3(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[73:37][3]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U4(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[73:37][4]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U5(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[73:37][5]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U6(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[73:37][6]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U7(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[73:37][7]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U8(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[73:37][8]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U9(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[73:37][9]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U10(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[73:37][10]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U11(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[73:37][11]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U12(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[73:37][12]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U13(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[73:37][13]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U14(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[73:37][14]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U15(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[73:37][15]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U16(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[73:37][16]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U17(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[73:37][17]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U18(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[73:37][18]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U19(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[73:37][19]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U20(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[73:37][20]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U21(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[73:37][21]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U22(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[73:37][22]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U23(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[73:37][23]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U24(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[73:37][24]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U25(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[73:37][25]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U26(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[73:37][26]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U27(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[73:37][27]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U28(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[73:37][28]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U29(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[73:37][29]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U30(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[73:37][30]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U31(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[73:37][31]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U32(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[73:37][32]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U33(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[73:37][33]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U34(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[73:37][34]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U35(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[73:37][35]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U36(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[73:37][36]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U321111(.IN1(int_req_v[73:37][0]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1 * 37)]), .S(and4resu_input_datapath1), .Q(int_req_v[73:37][0]));
	MUX21X1 U331112(.IN1(int_req_v[73:37][1]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+1]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+1]));
	MUX21X1 U331122(.IN1(int_req_v[73:37][2]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+2]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1]),.IN2(int_resp_v[2:1]), .S(and4resu_input_datapath1), .Q(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1+1]),.IN2(int_resp_v[2:1]), .S(and4resu_input_datapath1), .Q(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1+1]));

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule22[0]), .Y(next_read_ptr_fifomodule22[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule22[1]), .Y(next_read_ptr_fifomodule22[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule22[0]), .Y(next_write_ptr_fifomodule22[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule22[1]), .Y(next_write_ptr_fifomodule22[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule22[0]), .IN2(read_ptr_ff_fifomodule22[0]), .Q(u1temp_fifomodule22) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule22[1]), .IN2(read_ptr_ff_fifomodule22[1]), .Q(u2temp_fifomodule22) );
	AND2X1 U3 ( .A(u1temp_fifomodule22), .B(u2temp_fifomodule22), .Y(empty_vc_buffer22) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule22[1]), .B(read_ptr_ff_fifomodule22[1]), .Y(u4temp_fifomodule22) );
	AND2X1 U5 ( .A(u1temp_fifomodule22), .B(u4temp_fifomodule22), .Y(full_vc_buffer22) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][7]));

	INVX1 U7 ( .A(full_vc_buffer22), .Y(full_vc_buffer22_not_fifomodule) );
	AND2X1 U8 ( .A(write_flit22_vc_buffer2), .B(full_vc_buffer22_not_fifomodule), .Y(u7temp_fifomodule22) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule22), .Q(u9temp_fifomodule22));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule22[0]), .B0(u9temp_fifomodule22), .C1(u10carry_fifomodule22), .SO(next_write_ptr_fifomodule22[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule22), .B0(write_ptr_ff_fifomodule22[1]), .C1(u11carry_fifomodule22), .SO(next_write_ptr_fifomodule22[1]) );

	INVX1 U12 ( .A(empty_vc_buffer22), .Y(empty_vc_buffer22_not_fifomodule) );
	AND2X1 U13 ( .A(read_flit22_vc_buffer2), .B(empty_vc_buffer22_not_fifomodule), .Y(u13temp_fifomodule22) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule22), .Q(u14temp_fifomodule22));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule22[0]), .B0(u14temp_fifomodule22), .C1(u15carry_fifomodule22), .SO(next_read_ptr_fifomodule22[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule22), .B0(read_ptr_ff_fifomodule22[1]), .C1(u16carry_fifomodule22), .SO(next_read_ptr_fifomodule22[1]) );

	AND2X1 U17 ( .A(write_flit22_vc_buffer2), .B(full_vc_buffer22), .Y(u17res_fifomodule22) );
	AND2X1 U18 ( .A(read_flit22_vc_buffer2), .B(empty_vc_buffer22), .Y(u18res_fifomodule22) );
    OR2X1 U19 ( .A(u17res_fifomodule22), .B(u18res_fifomodule22), .Y(error_vc_buffer22) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule22[0]), .B(read_ptr_ff_fifomodule22[0]), .Y(fifo_ocup_fifomodule22[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule22[0]), .Y(write_ptr_ff_fifomodule22_0_not2) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule22_0_not2), .B(read_ptr_ff_fifomodule22[0]), .Y(b0wire_fifomodule22) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule22[1]), .B(read_ptr_ff_fifomodule22[1]), .Y(u23temp_fifomodule22) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule22[1]), .Y(write_ptr_ff_fifomodule22_1_not2) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule22[1]), .B(write_ptr_ff_fifomodule22_1_not2), .Y(boutb_fifomodule22) );
	XOR2X1 U24 ( .A(u23temp_fifomodule22), .B(b0wire_fifomodule22), .Y(fifo_ocup_fifomodule22[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule22), .Y(u23temp_fifomodule22_not_fifomodule22) );
	AND2X1 U26 ( .A(b0wire_fifomodule22), .B(u23temp_fifomodule22_not_fifomodule22), .Y(bouta_fifomodule22) );
	OR2X1 U27 ( .A(bouta_fifomodule22), .B(boutb_fifomodule22), .Y(boutmain_fifomodule22) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule22[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule22[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule22) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule22) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(write_ptr_ff_fifomodule22[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(read_ptr_ff_fifomodule22[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(fifo_ff_fifomodule22[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(write_ptr_ff_fifomodule22[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(read_ptr_ff_fifomodule22[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(fifo_ff_fifomodule22[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule22[0]), .Q(write_ptr_ff_fifomodule22[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule22[1]), .Q(write_ptr_ff_fifomodule22[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule22[0]), .Q(read_ptr_ff_fifomodule22[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule22[1]), .Q(read_ptr_ff_fifomodule22[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][0]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][1]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][2]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][3]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][4]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][5]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][6]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][7]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer22), .Y(next_locked_vc_buffer22) );
    BUFX1 U0(.A(flit22[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][0]));
	BUFX1 U1(.A(flit22[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][1]));
	BUFX1 U2(.A(flit22[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][2]));
	BUFX1 U3(.A(flit22[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][3]));
	BUFX1 U4(.A(flit22[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][4]));
	BUFX1 U5(.A(flit22[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][5]));
	BUFX1 U6(.A(flit22[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][6]));
	BUFX1 U7(.A(flit22[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][7]));
	BUFX1 U8(.A(flit22[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][8]));
	BUFX1 U9(.A(flit22[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][9]));
	BUFX1 U10(.A(flit22[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][10]));
	BUFX1 U11(.A(flit22[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][11]));
	BUFX1 U12(.A(flit22[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][12]));
	BUFX1 U13(.A(flit22[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][13]));
	BUFX1 U14(.A(flit22[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][14]));
	BUFX1 U15(.A(flit22[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][15]));
	BUFX1 U16(.A(flit22[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][16]));
	BUFX1 U17(.A(flit22[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][17]));
	BUFX1 U18(.A(flit22[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][18]));
	BUFX1 U19(.A(flit22[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][19]));
	BUFX1 U20(.A(flit22[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][20]));
	BUFX1 U21(.A(flit22[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][21]));
	BUFX1 U22(.A(flit22[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][22]));
	BUFX1 U23(.A(flit22[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][23]));
	BUFX1 U24(.A(flit22[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][24]));
	BUFX1 U25(.A(flit22[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][25]));
	BUFX1 U26(.A(flit22[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][26]));
	BUFX1 U27(.A(flit22[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][27]));
	BUFX1 U28(.A(flit22[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][28]));
	BUFX1 U29(.A(flit22[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][29]));
	BUFX1 U30(.A(flit22[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][30]));
	BUFX1 U31(.A(flit22[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][31]));
	BUFX1 U32(.A(flit22[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][32]));
	BUFX1 U33(.A(flit22[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][33]));
    NOR2X1 U34 ( .IN1(flit22[33]), .IN2(flit22[32]), .QN(norres_vc_buffer22_vc_buffer22) );
    OR4X1 U35 ( .IN1(flit22[29]), .IN2(flit22[28]), .IN3(flit22[27]), .IN4(flit22[26]), .Y(or1res_vc_buffer22) );
    OR4X1 U35 ( .IN1(flit22[25]), .IN2(flit22[24]), .IN3(flit22[23]), .IN4(flit22[22]), .Y(or2res_vc_buffer22) );
    OR2X1 U36 ( .A(or1res_vc_buffer22), .B(or2res_vc_buffer22), .Y(orres_vc_buffer22) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(norres_vc_buffer22_vc_buffer22), .IN3(orres_vc_buffer22), .Q(finres1_vc_buffer22) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer22), .IN2(1'b1), .S(finres1_vc_buffer22), .Q(next_locked_vc_buffer22);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(flit22[33]), .IN3(flit22[32]), .Q(andres1_vc_buffer22) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer22), .IN2(1'b0), .S(andres1_vc_buffer22), .Q(next_locked_vc_buffer22);

    INVX1 U41 ( .A(full_vc_buffer22), .Y(full_vc_buffer22_not) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer22), .Y(locked_by_route_ff_vc_buffer22_not) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer22_not), .S(norres_vc_buffer22_vc_buffer22), .Q(thirdand_vc_buffer22);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(full_vc_buffer22_not), .IN3(thirdand_vc_buffer22), .Q(write_flit22_vc_buffer2) );
    AND2X1 U45 ( .IN1(full_vc_buffer22_not), .IN2(norres_vc_buffer22_vc_buffer22), .Q(from_input_resp_input_datapath2[0]) );
    INVX1 U46 ( .A(empty_vc_buffer22), .Y(to_output_req_in_jump_input_datapath2put_datapath2[0]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[0]), .IN2(to_output_resp_input_datapath2[0]), .Q(read_flit22_vc_buffer2) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath2put_datapath2[2:1]), .Y(2'b00));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer22), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer22);

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule221[0]), .Y(next_read_ptr_fifomodule221[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule221[1]), .Y(next_read_ptr_fifomodule221[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule221[0]), .Y(next_write_ptr_fifomodule221[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule221[1]), .Y(next_write_ptr_fifomodule221[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule221[0]), .IN2(read_ptr_ff_fifomodule221[0]), .Q(u1temp_fifomodule221) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule221[1]), .IN2(read_ptr_ff_fifomodule221[1]), .Q(u2temp_fifomodule221) );
	AND2X1 U3 ( .A(u1temp_fifomodule221), .B(u2temp_fifomodule221), .Y(empty_vc_buffer221) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule221[1]), .B(read_ptr_ff_fifomodule221[1]), .Y(u4temp_fifomodule221) );
	AND2X1 U5 ( .A(u1temp_fifomodule221), .B(u4temp_fifomodule221), .Y(full_vc_buffer221) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][7]));

	INVX1 U7 ( .A(full_vc_buffer221), .Y(full_vc_buffer221_not1_fifomodule1) );
	AND2X1 U8 ( .A(write_flit221_vc_buffer12), .B(full_vc_buffer221_not1_fifomodule1), .Y(u7temp_fifomodule221) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule221), .Q(u9temp_fifomodule221));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule221[0]), .B0(u9temp_fifomodule221), .C1(u10carry_fifomodule221), .SO(next_write_ptr_fifomodule221[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule221), .B0(write_ptr_ff_fifomodule221[1]), .C1(u11carry_fifomodule221), .SO(next_write_ptr_fifomodule221[1]) );

	INVX1 U12 ( .A(empty_vc_buffer221), .Y(empty_vc_buffer221_not_fifomodule1) );
	AND2X1 U13 ( .A(read_flit221_vc_buffer12), .B(empty_vc_buffer221_not_fifomodule1), .Y(u13temp_fifomodule221) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule221), .Q(u14temp_fifomodule221));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule221[0]), .B0(u14temp_fifomodule221), .C1(u15carry_fifomodule221), .SO(next_read_ptr_fifomodule221[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule221), .B0(read_ptr_ff_fifomodule221[1]), .C1(u16carry_fifomodule221), .SO(next_read_ptr_fifomodule221[1]) );

	AND2X1 U17 ( .A(write_flit221_vc_buffer12), .B(full_vc_buffer221), .Y(u17res_fifomodule221) );
	AND2X1 U18 ( .A(read_flit221_vc_buffer12), .B(empty_vc_buffer221), .Y(u18res_fifomodule221) );
    OR2X1 U19 ( .A(u17res_fifomodule221), .B(u18res_fifomodule221), .Y(error_vc_buffer221) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule221[0]), .B(read_ptr_ff_fifomodule221[0]), .Y(fifo_ocup_fifomodule221[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule221[0]), .Y(write_ptr_ff_fifomodule221_0_not12) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule221_0_not12), .B(read_ptr_ff_fifomodule221[0]), .Y(b0wire_fifomodule221) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule221[1]), .B(read_ptr_ff_fifomodule221[1]), .Y(u23temp_fifomodule221) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule221[1]), .Y(write_ptr_ff_fifomodule221_1_not12) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule221[1]), .B(write_ptr_ff_fifomodule221_1_not12), .Y(boutb_fifomodule221) );
	XOR2X1 U24 ( .A(u23temp_fifomodule221), .B(b0wire_fifomodule221), .Y(fifo_ocup_fifomodule221[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule221), .Y(u23temp_fifomodule221_not_fifomodule1) );
	AND2X1 U26 ( .A(b0wire_fifomodule221), .B(u23temp_fifomodule221_not_fifomodule1), .Y(bouta_fifomodule221) );
	OR2X1 U27 ( .A(bouta_fifomodule221), .B(boutb_fifomodule221), .Y(boutmain_fifomodule221) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule221[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule221[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule221) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule221) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(write_ptr_ff_fifomodule221[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(read_ptr_ff_fifomodule221[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(fifo_ff_fifomodule221[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(write_ptr_ff_fifomodule221[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(read_ptr_ff_fifomodule221[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(fifo_ff_fifomodule221[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule221[0]), .Q(write_ptr_ff_fifomodule221[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule221[1]), .Q(write_ptr_ff_fifomodule221[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule221[0]), .Q(read_ptr_ff_fifomodule221[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule221[1]), .Q(read_ptr_ff_fifomodule221[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][0]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][1]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][2]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][3]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][4]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][5]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][6]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][7]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer221), .Y(next_locked_vc_buffer221) );
    BUFX1 U0(.A(flit221[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][0]));
	BUFX1 U1(.A(flit221[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][1]));
	BUFX1 U2(.A(flit221[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][2]));
	BUFX1 U3(.A(flit221[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][3]));
	BUFX1 U4(.A(flit221[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][4]));
	BUFX1 U5(.A(flit221[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][5]));
	BUFX1 U6(.A(flit221[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][6]));
	BUFX1 U7(.A(flit221[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][7]));
	BUFX1 U8(.A(flit221[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][8]));
	BUFX1 U9(.A(flit221[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][9]));
	BUFX1 U10(.A(flit221[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][10]));
	BUFX1 U11(.A(flit221[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][11]));
	BUFX1 U12(.A(flit221[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][12]));
	BUFX1 U13(.A(flit221[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][13]));
	BUFX1 U14(.A(flit221[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][14]));
	BUFX1 U15(.A(flit221[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][15]));
	BUFX1 U16(.A(flit221[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][16]));
	BUFX1 U17(.A(flit221[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][17]));
	BUFX1 U18(.A(flit221[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][18]));
	BUFX1 U19(.A(flit221[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][19]));
	BUFX1 U20(.A(flit221[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][20]));
	BUFX1 U21(.A(flit221[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][21]));
	BUFX1 U22(.A(flit221[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][22]));
	BUFX1 U23(.A(flit221[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][23]));
	BUFX1 U24(.A(flit221[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][24]));
	BUFX1 U25(.A(flit221[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][25]));
	BUFX1 U26(.A(flit221[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][26]));
	BUFX1 U27(.A(flit221[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][27]));
	BUFX1 U28(.A(flit221[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][28]));
	BUFX1 U29(.A(flit221[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][29]));
	BUFX1 U30(.A(flit221[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][30]));
	BUFX1 U31(.A(flit221[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][31]));
	BUFX1 U32(.A(flit221[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][32]));
	BUFX1 U33(.A(flit221[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][33]));
    NOR2X1 U34 ( .IN1(flit221[33]), .IN2(flit221[32]), .QN(norres_vc_buffer221_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit221[29]), .IN2(flit221[28]), .IN3(flit221[27]), .IN4(flit221[26]), .Y(or1res_vc_buffer221) );
    OR4X1 U35 ( .IN1(flit221[25]), .IN2(flit221[24]), .IN3(flit221[23]), .IN4(flit221[22]), .Y(or2res_vc_buffer221) );
    OR2X1 U36 ( .A(or1res_vc_buffer221), .B(or2res_vc_buffer221), .Y(orres_vc_buffer221) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(norres_vc_buffer221_vc_buffer1), .IN3(orres_vc_buffer221), .Q(finres1_vc_buffer221) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer221), .IN2(1'b1), .S(finres1_vc_buffer221), .Q(next_locked_vc_buffer221);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(flit221[33]), .IN3(flit221[32]), .Q(andres1_vc_buffer221) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer221), .IN2(1'b0), .S(andres1_vc_buffer221), .Q(next_locked_vc_buffer221);

    INVX1 U41 ( .A(full_vc_buffer221), .Y(full_vc_buffer221_not1) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer221), .Y(locked_by_route_ff_vc_buffer221_not1) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer221_not1), .S(norres_vc_buffer221_vc_buffer1), .Q(thirdand_vc_buffer221);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(full_vc_buffer221_not1), .IN3(thirdand_vc_buffer221), .Q(write_flit221_vc_buffer12) );
    AND2X1 U45 ( .IN1(full_vc_buffer221_not1), .IN2(norres_vc_buffer221_vc_buffer1), .Q(from_input_resp_input_datapath2[1]) );
    INVX1 U46 ( .A(empty_vc_buffer221), .Y(to_output_req_in_jump_input_datapath2put_datapath2[37]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[37]), .IN2(to_output_resp_input_datapath2[1]), .Q(read_flit221_vc_buffer12) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath2put_datapath2[39:38]), .Y(2'b01));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer221), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer221);


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule222[0]), .Y(next_read_ptr_fifomodule222[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule222[1]), .Y(next_read_ptr_fifomodule222[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule222[0]), .Y(next_write_ptr_fifomodule222[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule222[1]), .Y(next_write_ptr_fifomodule222[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule222[0]), .IN2(read_ptr_ff_fifomodule222[0]), .Q(u1temp_fifomodule222) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule222[1]), .IN2(read_ptr_ff_fifomodule222[1]), .Q(u2temp_fifomodule222) );
	AND2X1 U3 ( .A(u1temp_fifomodule222), .B(u2temp_fifomodule222), .Y(empty_vc_buffer222) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule222[1]), .B(read_ptr_ff_fifomodule222[1]), .Y(u4temp_fifomodule222) );
	AND2X1 U5 ( .A(u1temp_fifomodule222), .B(u4temp_fifomodule222), .Y(full_vc_buffer222) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][7]));

	INVX1 U7 ( .A(full_vc_buffer222), .Y(full_vc_buffer222_not2_fifomodule2) );
	AND2X1 U8 ( .A(write_flit222_vc_buffer22), .B(full_vc_buffer222_not2_fifomodule2), .Y(u7temp_fifomodule222) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule222), .Q(u9temp_fifomodule222));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule222[0]), .B0(u9temp_fifomodule222), .C1(u10carry_fifomodule222), .SO(next_write_ptr_fifomodule222[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule222), .B0(write_ptr_ff_fifomodule222[1]), .C1(u11carry_fifomodule222), .SO(next_write_ptr_fifomodule222[1]) );

	INVX1 U12 ( .A(empty_vc_buffer222), .Y(empty_vc_buffer222_not_fifomodule2) );
	AND2X1 U13 ( .A(read_flit222_vc_buffer22), .B(empty_vc_buffer222_not_fifomodule2), .Y(u13temp_fifomodule222) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule222), .Q(u14temp_fifomodule222));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule222[0]), .B0(u14temp_fifomodule222), .C1(u15carry_fifomodule222), .SO(next_read_ptr_fifomodule222[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule222), .B0(read_ptr_ff_fifomodule222[1]), .C1(u16carry_fifomodule222), .SO(next_read_ptr_fifomodule222[1]) );

	AND2X1 U17 ( .A(write_flit222_vc_buffer22), .B(full_vc_buffer222), .Y(u17res_fifomodule222) );
	AND2X1 U18 ( .A(read_flit222_vc_buffer22), .B(empty_vc_buffer222), .Y(u18res_fifomodule222) );
    OR2X1 U19 ( .A(u17res_fifomodule222), .B(u18res_fifomodule222), .Y(error_vc_buffer222) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule222[0]), .B(read_ptr_ff_fifomodule222[0]), .Y(fifo_ocup_fifomodule222[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule222[0]), .Y(write_ptr_ff_fifomodule222_0_not22) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule222_0_not22), .B(read_ptr_ff_fifomodule222[0]), .Y(b0wire_fifomodule222) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule222[1]), .B(read_ptr_ff_fifomodule222[1]), .Y(u23temp_fifomodule222) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule222[1]), .Y(write_ptr_ff_fifomodule222_1_not22) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule222[1]), .B(write_ptr_ff_fifomodule222_1_not22), .Y(boutb_fifomodule222) );
	XOR2X1 U24 ( .A(u23temp_fifomodule222), .B(b0wire_fifomodule222), .Y(fifo_ocup_fifomodule222[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule222), .Y(u23temp_fifomodule222_not_fifomodule2) );
	AND2X1 U26 ( .A(b0wire_fifomodule222), .B(u23temp_fifomodule222_not_fifomodule2), .Y(bouta_fifomodule222) );
	OR2X1 U27 ( .A(bouta_fifomodule222), .B(boutb_fifomodule222), .Y(boutmain_fifomodule222) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule222[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule222[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule222) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule222) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(write_ptr_ff_fifomodule222[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(read_ptr_ff_fifomodule222[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(fifo_ff_fifomodule222[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(write_ptr_ff_fifomodule222[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(read_ptr_ff_fifomodule222[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(fifo_ff_fifomodule222[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule222[0]), .Q(write_ptr_ff_fifomodule222[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule222[1]), .Q(write_ptr_ff_fifomodule222[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule222[0]), .Q(read_ptr_ff_fifomodule222[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule222[1]), .Q(read_ptr_ff_fifomodule222[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][0]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][1]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][2]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][3]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][4]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][5]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][6]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][7]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer222), .Y(next_locked_vc_buffer222) );
    BUFX1 U0(.A(flit222[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][0]));
	BUFX1 U1(.A(flit222[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][1]));
	BUFX1 U2(.A(flit222[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][2]));
	BUFX1 U3(.A(flit222[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][3]));
	BUFX1 U4(.A(flit222[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][4]));
	BUFX1 U5(.A(flit222[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][5]));
	BUFX1 U6(.A(flit222[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][6]));
	BUFX1 U7(.A(flit222[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][7]));
	BUFX1 U8(.A(flit222[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][8]));
	BUFX1 U9(.A(flit222[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][9]));
	BUFX1 U10(.A(flit222[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][10]));
	BUFX1 U11(.A(flit222[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][11]));
	BUFX1 U12(.A(flit222[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][12]));
	BUFX1 U13(.A(flit222[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][13]));
	BUFX1 U14(.A(flit222[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][14]));
	BUFX1 U15(.A(flit222[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][15]));
	BUFX1 U16(.A(flit222[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][16]));
	BUFX1 U17(.A(flit222[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][17]));
	BUFX1 U18(.A(flit222[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][18]));
	BUFX1 U19(.A(flit222[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][19]));
	BUFX1 U20(.A(flit222[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][20]));
	BUFX1 U21(.A(flit222[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][21]));
	BUFX1 U22(.A(flit222[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][22]));
	BUFX1 U23(.A(flit222[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][23]));
	BUFX1 U24(.A(flit222[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][24]));
	BUFX1 U25(.A(flit222[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][25]));
	BUFX1 U26(.A(flit222[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][26]));
	BUFX1 U27(.A(flit222[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][27]));
	BUFX1 U28(.A(flit222[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][28]));
	BUFX1 U29(.A(flit222[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][29]));
	BUFX1 U30(.A(flit222[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][30]));
	BUFX1 U31(.A(flit222[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][31]));
	BUFX1 U32(.A(flit222[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][32]));
	BUFX1 U33(.A(flit222[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][33]));
    NOR2X1 U34 ( .IN1(flit222[33]), .IN2(flit222[32]), .QN(norres_vc_buffer222_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit222[29]), .IN2(flit222[28]), .IN3(flit222[27]), .IN4(flit222[26]), .Y(or1res_vc_buffer222) );
    OR4X1 U35 ( .IN1(flit222[25]), .IN2(flit222[24]), .IN3(flit222[23]), .IN4(flit222[22]), .Y(or2res_vc_buffer222) );
    OR2X1 U36 ( .A(or1res_vc_buffer222), .B(or2res_vc_buffer222), .Y(orres_vc_buffer222) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(norres_vc_buffer222_vc_buffer2), .IN3(orres_vc_buffer222), .Q(finres1_vc_buffer222) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer222), .IN2(1'b1), .S(finres1_vc_buffer222), .Q(next_locked_vc_buffer222);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(flit222[33]), .IN3(flit222[32]), .Q(andres1_vc_buffer222) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer222), .IN2(1'b0), .S(andres1_vc_buffer222), .Q(next_locked_vc_buffer222);

    INVX1 U41 ( .A(full_vc_buffer222), .Y(full_vc_buffer222_not2) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer222), .Y(locked_by_route_ff_vc_buffer222_not2) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer222_not2), .S(norres_vc_buffer222_vc_buffer2), .Q(thirdand_vc_buffer222);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(full_vc_buffer222_not2), .IN3(thirdand_vc_buffer222), .Q(write_flit222_vc_buffer22) );
    AND2X1 U45 ( .IN1(full_vc_buffer222_not2), .IN2(norres_vc_buffer222_vc_buffer2), .Q(from_input_resp_input_datapath2[2]) );
    INVX1 U46 ( .A(empty_vc_buffer222), .Y(to_output_req_in_jump_input_datapath2put_datapath2[74]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[74]), .IN2(to_output_resp_input_datapath2[2]), .Q(read_flit222_vc_buffer22) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath2put_datapath2[76:75]), .Y(2'b10));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer222), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer222);

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath2put_datapath2[77]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath2put_datapath2[78]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath2put_datapath2[79]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath2put_datapath2[80]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath2put_datapath2[81]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath2put_datapath2[82]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath2put_datapath2[83]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath2put_datapath2[84]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath2put_datapath2[85]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath2put_datapath2[86]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath2put_datapath2[87]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath2put_datapath2[88]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath2put_datapath2[89]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath2put_datapath2[90]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath2put_datapath2[91]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath2put_datapath2[92]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath2put_datapath2[93]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath2put_datapath2[94]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath2put_datapath2[95]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath2put_datapath2[96]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath2put_datapath2[97]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath2put_datapath2[98]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath2put_datapath2[99]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath2put_datapath2[100]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath2put_datapath2[101]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath2put_datapath2[102]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath2put_datapath2[103]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath2put_datapath2[104]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath2put_datapath2[105]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath2put_datapath2[106]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath2put_datapath2[107]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath2put_datapath2[108]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath2put_datapath2[109]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath2put_datapath2[110]), .Y(ext_req_v_i[110:74][36]));
    XNOR2X1 U222 ( .IN1(ext_req_v_i[110:74][1]), .IN2(i_input_datapath2[0]), .QN(xnor1resu_input_datapath2) );
    XNOR2X1 U222 ( .IN1(ext_req_v_i[110:74][2]), .IN2(i_input_datapath2[1]), .QN(xnor2resu_input_datapath2) );
    AND2X1 U128 ( .IN1(xnor1resu_input_datapath2), .IN2(xnor2resu_input_datapath2), .Q(and1resu_input_datapath2) );
    AND3X1 U128 ( .IN1(and1resu_input_datapath2), .IN2(ext_req_v_i[110:74][0]), .IN2(ext_req_v_i[110:74][0]), .Q(cond1line_input_datapath2) );
    MUX21X1 U0009 (.IN1(vc_ch_act_in_input_datapath2[0]), .IN2(i_input_datapath2[0]), .S(cond1line_input_datapath2), .Q(vc_ch_act_in_input_datapath2[0]));
    MUX21X1 U0010 (.IN1(vc_ch_act_in_input_datapath2[1]), .IN2(i_input_datapath2[1]), .S(cond1line_input_datapath2), .Q(vc_ch_act_in_input_datapath2[1]));
    MUX21X1 U0011 (.IN1(req_in_jump_input_datapath2), .IN2(1), .S(cond1line_input_datapath2), .Q(req_in_jump_input_datapath2));
	BUFX1 U3(.A(from_input_req_in_jump_input_datapath2put_datapath2[40]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath2put_datapath2[41]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath2put_datapath2[42]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath2put_datapath2[43]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath2put_datapath2[44]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath2put_datapath2[45]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath2put_datapath2[46]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath2put_datapath2[47]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath2put_datapath2[48]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath2put_datapath2[49]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath2put_datapath2[50]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath2put_datapath2[51]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath2put_datapath2[52]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath2put_datapath2[53]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath2put_datapath2[54]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath2put_datapath2[55]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath2put_datapath2[56]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath2put_datapath2[57]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath2put_datapath2[58]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath2put_datapath2[59]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath2put_datapath2[60]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath2put_datapath2[61]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath2put_datapath2[62]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath2put_datapath2[63]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath2put_datapath2[64]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath2put_datapath2[65]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath2put_datapath2[66]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath2put_datapath2[67]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath2put_datapath2[68]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath2put_datapath2[69]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath2put_datapath2[70]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath2put_datapath2[71]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath2put_datapath2[72]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath2put_datapath2[73]), .Y(ext_req_v_i[110:74][36]));

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath2put_datapath2[3]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath2put_datapath2[4]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath2put_datapath2[5]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath2put_datapath2[6]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath2put_datapath2[7]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath2put_datapath2[8]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath2put_datapath2[9]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath2put_datapath2[10]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath2put_datapath2[11]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath2put_datapath2[12]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath2put_datapath2[13]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath2put_datapath2[14]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath2put_datapath2[15]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath2put_datapath2[16]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath2put_datapath2[17]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath2put_datapath2[18]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath2put_datapath2[19]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath2put_datapath2[20]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath2put_datapath2[21]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath2put_datapath2[22]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath2put_datapath2[23]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath2put_datapath2[24]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath2put_datapath2[25]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath2put_datapath2[26]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath2put_datapath2[27]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath2put_datapath2[28]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath2put_datapath2[29]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath2put_datapath2[30]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath2put_datapath2[31]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath2put_datapath2[32]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath2put_datapath2[33]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath2put_datapath2[34]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath2put_datapath2[35]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath2put_datapath2[36]), .Y(ext_req_v_i[110:74][36]));

    MUX21X1 U0012 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2 * 37]), .IN2(ext_req_v_i[110:74][0]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2 * 37]));
    MUX21X1 U0013 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+2]), .IN2(vc_ch_act_in_input_datapath2[1]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+2]));
    MUX21X1 U0014 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+1]), .IN2(vc_ch_act_in_input_datapath2[0]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+1]));
    MUX21X1 U0015 (.IN1(ext_resp_v_o[3:2][0]), .IN2(from_input_resp_input_datapath2[vc_ch_act_in_input_datapath2]), .S(req_in_jump_input_datapath2), .Q(ext_resp_v_o[3:2][0]));

    INVX1 U041 ( .A(req_in_jump_input_datapath2), .Y(req_in_jump_input_datapath2_not) );
    MUX21X1 U0016 (.IN1(ext_resp_v_o[3:2][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath2_not), .Q(ext_resp_v_o[3:2][0]));
    BUFX1 U34(.A(from_input_req_in_jump_input_datapath2put_datapath2[34]), .Y(ext_req_v_i[110:74][34]));

    XOR2X1 U0222 ( .IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b1), .Q(xor1resu_input_datapath2) );
    MUX21X1 U0017 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(xor1resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U0018 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b0), .S(xor1resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[1]));
    AND2X1 U38123 ( .IN1(xor1resu_input_datapath2), .IN2(to_output_req_in_jump_input_datapath2put_datapath2[j_input_datapath2*37]), .Q(and2resu_input_datapath2) );
    MUX21X1 U0019 (.IN1(vc_ch_act_out_input_datapath2[0]), .IN2(j_input_datapath2[0]), .S(and2resu_input_datapath2), .Q(vc_ch_act_out_input_datapath2[0]));
    MUX21X1 U0020 (.IN1(vc_ch_act_out_input_datapath2[1]), .IN2(j_input_datapath2[1]), .S(and2resu_input_datapath2), .Q(vc_ch_act_out_input_datapath2[1]));
    MUX21X1 U0021 (.IN1(req_out_jump_input_datapath2), .IN2(1'b1), .S(and2resu_input_datapath2), .Q(req_out_jump_input_datapath2));
    MUX21X1 U0022 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(and2resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U0023 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b1), .S(and2resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[1]));
    HADDX1 U00021 ( .A0(j_input_datapath2[0]), .B0(1'b1), .C1(j_input_datapath2[1]), .SO(j_input_datapath2[0]) );
    HADDX1 U00022 ( .A0(j_input_datapath2[0]), .B0(1'b1), .C1(j_input_datapath2[1]), .SO(j_input_datapath2[0]) );
    AND2X1 U38111 ( .IN1(xor1resu_input_datapath2), .IN2(to_output_req_in_jump_input_datapath2put_datapath2[j_input_datapath2*37]), .Q(and3resu) );
    NAND2X1 U29311(.A(_sv2v_jump_input_datapath2[0]),.B(_sv2v_jump_input_datapath2[1]),.Y(nand1resu_input_datapath22));
    MUX21X1 U00212 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(nand1resu_input_datapath22), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U00213 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b0), .S(nand1resu_input_datapath22), .Q(_sv2v_jump_input_datapath2[1]));
    XNOR2X1 U17581 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(_sv2v_jump_input_datapath2[1]), .Q(xnor23resu_input_datapath2) );
    AND2X1 U38111 ( .IN1(xnor23resu_input_datapath2), .IN2(req_out_jump_input_datapath2), .Q(and4resu_input_datapath2) );

    MUX21X1 U3(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[110:74][3]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U4(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[110:74][4]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U5(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[110:74][5]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U6(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[110:74][6]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U7(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[110:74][7]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U8(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[110:74][8]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U9(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[110:74][9]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U10(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[110:74][10]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U11(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[110:74][11]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U12(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[110:74][12]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U13(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[110:74][13]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U14(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[110:74][14]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U15(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[110:74][15]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U16(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[110:74][16]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U17(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[110:74][17]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U18(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[110:74][18]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U19(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[110:74][19]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U20(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[110:74][20]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U21(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[110:74][21]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U22(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[110:74][22]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U23(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[110:74][23]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U24(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[110:74][24]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U25(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[110:74][25]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U26(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[110:74][26]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U27(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[110:74][27]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U28(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[110:74][28]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U29(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[110:74][29]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U30(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[110:74][30]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U31(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[110:74][31]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U32(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[110:74][32]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U33(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[110:74][33]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U34(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[110:74][34]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U35(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[110:74][35]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U36(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[110:74][36]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U321111(.IN1(int_req_v[110:74][0]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2 * 37)]), .S(and4resu_input_datapath2), .Q(int_req_v[110:74][0]));
	MUX21X1 U331112(.IN1(int_req_v[110:74][1]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+1]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+1]));
	MUX21X1 U331122(.IN1(int_req_v[110:74][2]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+2]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2]),.IN2(int_resp_v[3:2]), .S(and4resu_input_datapath2), .Q(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2+1]),.IN2(int_resp_v[3:2]), .S(and4resu_input_datapath2), .Q(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2+1]));


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule3[0]), .Y(next_read_ptr_fifomodule3[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule3[1]), .Y(next_read_ptr_fifomodule3[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule3[0]), .Y(next_write_ptr_fifomodule3[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule3[1]), .Y(next_write_ptr_fifomodule3[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule3[0]), .IN2(read_ptr_ff_fifomodule3[0]), .Q(u1temp_fifomodule3) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule3[1]), .IN2(read_ptr_ff_fifomodule3[1]), .Q(u2temp_fifomodule3) );
	AND2X1 U3 ( .A(u1temp_fifomodule3), .B(u2temp_fifomodule3), .Y(empty_vc_buffer3) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule3[1]), .B(read_ptr_ff_fifomodule3[1]), .Y(u4temp_fifomodule3) );
	AND2X1 U5 ( .A(u1temp_fifomodule3), .B(u4temp_fifomodule3), .Y(full_vc_buffer3) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][7]));

	INVX1 U7 ( .A(full_vc_buffer3), .Y(full_vc_buffer3_not_fifomodule) );
	AND2X1 U8 ( .A(write_flit3_vc_buffer3), .B(full_vc_buffer3_not_fifomodule), .Y(u7temp_fifomodule3) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule3), .Q(u9temp_fifomodule3));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule3[0]), .B0(u9temp_fifomodule3), .C1(u10carry_fifomodule3), .SO(next_write_ptr_fifomodule3[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule3), .B0(write_ptr_ff_fifomodule3[1]), .C1(u11carry_fifomodule3), .SO(next_write_ptr_fifomodule3[1]) );

	INVX1 U12 ( .A(empty_vc_buffer3), .Y(empty_vc_buffer3_not_fifomodule) );
	AND2X1 U13 ( .A(read_flit3_vc_buffer3), .B(empty_vc_buffer3_not_fifomodule), .Y(u13temp_fifomodule3) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule3), .Q(u14temp_fifomodule3));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule3[0]), .B0(u14temp_fifomodule3), .C1(u15carry_fifomodule3), .SO(next_read_ptr_fifomodule3[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule3), .B0(read_ptr_ff_fifomodule3[1]), .C1(u16carry_fifomodule3), .SO(next_read_ptr_fifomodule3[1]) );

	AND2X1 U17 ( .A(write_flit3_vc_buffer3), .B(full_vc_buffer3), .Y(u17res_fifomodule3) );
	AND2X1 U18 ( .A(read_flit3_vc_buffer3), .B(empty_vc_buffer3), .Y(u18res_fifomodule3) );
    OR2X1 U19 ( .A(u17res_fifomodule3), .B(u18res_fifomodule3), .Y(error_vc_buffer3) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule3[0]), .B(read_ptr_ff_fifomodule3[0]), .Y(fifo_ocup_fifomodule3[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule3[0]), .Y(write_ptr_ff_fifomodule3_0_not3) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule3_0_not3), .B(read_ptr_ff_fifomodule3[0]), .Y(b0wire_fifomodule3) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule3[1]), .B(read_ptr_ff_fifomodule3[1]), .Y(u23temp_fifomodule3) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule3[1]), .Y(write_ptr_ff_fifomodule3_1_not3) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule3[1]), .B(write_ptr_ff_fifomodule3_1_not3), .Y(boutb_fifomodule3) );
	XOR2X1 U24 ( .A(u23temp_fifomodule3), .B(b0wire_fifomodule3), .Y(fifo_ocup_fifomodule3[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule3), .Y(u23temp_fifomodule3_not_fifomodule3) );
	AND2X1 U26 ( .A(b0wire_fifomodule3), .B(u23temp_fifomodule3_not_fifomodule3), .Y(bouta_fifomodule3) );
	OR2X1 U27 ( .A(bouta_fifomodule3), .B(boutb_fifomodule3), .Y(boutmain_fifomodule3) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule3[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule3[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule3) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule3) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(write_ptr_ff_fifomodule3[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(read_ptr_ff_fifomodule3[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(fifo_ff_fifomodule3[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(write_ptr_ff_fifomodule3[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(read_ptr_ff_fifomodule3[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(fifo_ff_fifomodule3[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule3[0]), .Q(write_ptr_ff_fifomodule3[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule3[1]), .Q(write_ptr_ff_fifomodule3[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule3[0]), .Q(read_ptr_ff_fifomodule3[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule3[1]), .Q(read_ptr_ff_fifomodule3[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][0]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][1]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][2]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][3]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][4]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][5]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][6]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][7]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer3), .Y(next_locked_vc_buffer3) );
    BUFX1 U0(.A(flit3[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][0]));
	BUFX1 U1(.A(flit3[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][1]));
	BUFX1 U2(.A(flit3[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][2]));
	BUFX1 U3(.A(flit3[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][3]));
	BUFX1 U4(.A(flit3[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][4]));
	BUFX1 U5(.A(flit3[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][5]));
	BUFX1 U6(.A(flit3[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][6]));
	BUFX1 U7(.A(flit3[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][7]));
	BUFX1 U8(.A(flit3[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][8]));
	BUFX1 U9(.A(flit3[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][9]));
	BUFX1 U10(.A(flit3[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][10]));
	BUFX1 U11(.A(flit3[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][11]));
	BUFX1 U12(.A(flit3[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][12]));
	BUFX1 U13(.A(flit3[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][13]));
	BUFX1 U14(.A(flit3[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][14]));
	BUFX1 U15(.A(flit3[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][15]));
	BUFX1 U16(.A(flit3[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][16]));
	BUFX1 U17(.A(flit3[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][17]));
	BUFX1 U18(.A(flit3[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][18]));
	BUFX1 U19(.A(flit3[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][19]));
	BUFX1 U20(.A(flit3[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][20]));
	BUFX1 U21(.A(flit3[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][21]));
	BUFX1 U22(.A(flit3[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][22]));
	BUFX1 U23(.A(flit3[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][23]));
	BUFX1 U24(.A(flit3[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][24]));
	BUFX1 U25(.A(flit3[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][25]));
	BUFX1 U26(.A(flit3[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][26]));
	BUFX1 U27(.A(flit3[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][27]));
	BUFX1 U28(.A(flit3[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][28]));
	BUFX1 U29(.A(flit3[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][29]));
	BUFX1 U30(.A(flit3[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][30]));
	BUFX1 U31(.A(flit3[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][31]));
	BUFX1 U32(.A(flit3[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][32]));
	BUFX1 U33(.A(flit3[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][33]));
    NOR2X1 U34 ( .IN1(flit3[33]), .IN2(flit3[32]), .QN(norres_vc_buffer3_vc_buffer3) );
    OR4X1 U35 ( .IN1(flit3[29]), .IN2(flit3[28]), .IN3(flit3[27]), .IN4(flit3[26]), .Y(or1res_vc_buffer3) );
    OR4X1 U35 ( .IN1(flit3[25]), .IN2(flit3[24]), .IN3(flit3[23]), .IN4(flit3[22]), .Y(or2res_vc_buffer3) );
    OR2X1 U36 ( .A(or1res_vc_buffer3), .B(or2res_vc_buffer3), .Y(orres_vc_buffer3) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(norres_vc_buffer3_vc_buffer3), .IN3(orres_vc_buffer3), .Q(finres1_vc_buffer3) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer3), .IN2(1'b1), .S(finres1_vc_buffer3), .Q(next_locked_vc_buffer3);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(flit3[33]), .IN3(flit3[32]), .Q(andres1_vc_buffer3) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer3), .IN2(1'b0), .S(andres1_vc_buffer3), .Q(next_locked_vc_buffer3);

    INVX1 U41 ( .A(full_vc_buffer3), .Y(full_vc_buffer3_not) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer3), .Y(locked_by_route_ff_vc_buffer3_not) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer3_not), .S(norres_vc_buffer3_vc_buffer3), .Q(thirdand_vc_buffer3);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(full_vc_buffer3_not), .IN3(thirdand_vc_buffer3), .Q(write_flit3_vc_buffer3) );
    AND2X1 U45 ( .IN1(full_vc_buffer3_not), .IN2(norres_vc_buffer3_vc_buffer3), .Q(from_input_resp_input_datapath3[0]) );
    INVX1 U46 ( .A(empty_vc_buffer3), .Y(to_output_req_in_jump_input_datapath3put_datapath3[0]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[0]), .IN2(to_output_resp_input_datapath3[0]), .Q(read_flit3_vc_buffer3) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath3put_datapath3[2:1]), .Y(2'b00));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer3), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer3);

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule31[0]), .Y(next_read_ptr_fifomodule31[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule31[1]), .Y(next_read_ptr_fifomodule31[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule31[0]), .Y(next_write_ptr_fifomodule31[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule31[1]), .Y(next_write_ptr_fifomodule31[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule31[0]), .IN2(read_ptr_ff_fifomodule31[0]), .Q(u1temp_fifomodule31) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule31[1]), .IN2(read_ptr_ff_fifomodule31[1]), .Q(u2temp_fifomodule31) );
	AND2X1 U3 ( .A(u1temp_fifomodule31), .B(u2temp_fifomodule31), .Y(empty_vc_buffer31) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule31[1]), .B(read_ptr_ff_fifomodule31[1]), .Y(u4temp_fifomodule31) );
	AND2X1 U5 ( .A(u1temp_fifomodule31), .B(u4temp_fifomodule31), .Y(full_vc_buffer31) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][7]));

	INVX1 U7 ( .A(full_vc_buffer31), .Y(full_vc_buffer31_not1_fifomodule1) );
	AND2X1 U8 ( .A(write_flit31_vc_buffer13), .B(full_vc_buffer31_not1_fifomodule1), .Y(u7temp_fifomodule31) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule31), .Q(u9temp_fifomodule31));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule31[0]), .B0(u9temp_fifomodule31), .C1(u10carry_fifomodule31), .SO(next_write_ptr_fifomodule31[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule31), .B0(write_ptr_ff_fifomodule31[1]), .C1(u11carry_fifomodule31), .SO(next_write_ptr_fifomodule31[1]) );

	INVX1 U12 ( .A(empty_vc_buffer31), .Y(empty_vc_buffer31_not_fifomodule1) );
	AND2X1 U13 ( .A(read_flit31_vc_buffer13), .B(empty_vc_buffer31_not_fifomodule1), .Y(u13temp_fifomodule31) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule31), .Q(u14temp_fifomodule31));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule31[0]), .B0(u14temp_fifomodule31), .C1(u15carry_fifomodule31), .SO(next_read_ptr_fifomodule31[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule31), .B0(read_ptr_ff_fifomodule31[1]), .C1(u16carry_fifomodule31), .SO(next_read_ptr_fifomodule31[1]) );

	AND2X1 U17 ( .A(write_flit31_vc_buffer13), .B(full_vc_buffer31), .Y(u17res_fifomodule31) );
	AND2X1 U18 ( .A(read_flit31_vc_buffer13), .B(empty_vc_buffer31), .Y(u18res_fifomodule31) );
    OR2X1 U19 ( .A(u17res_fifomodule31), .B(u18res_fifomodule31), .Y(error_vc_buffer31) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule31[0]), .B(read_ptr_ff_fifomodule31[0]), .Y(fifo_ocup_fifomodule31[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule31[0]), .Y(write_ptr_ff_fifomodule31_0_not13) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule31_0_not13), .B(read_ptr_ff_fifomodule31[0]), .Y(b0wire_fifomodule31) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule31[1]), .B(read_ptr_ff_fifomodule31[1]), .Y(u23temp_fifomodule31) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule31[1]), .Y(write_ptr_ff_fifomodule31_1_not13) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule31[1]), .B(write_ptr_ff_fifomodule31_1_not13), .Y(boutb_fifomodule31) );
	XOR2X1 U24 ( .A(u23temp_fifomodule31), .B(b0wire_fifomodule31), .Y(fifo_ocup_fifomodule31[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule31), .Y(u23temp_fifomodule31_not_fifomodule1) );
	AND2X1 U26 ( .A(b0wire_fifomodule31), .B(u23temp_fifomodule31_not_fifomodule1), .Y(bouta_fifomodule31) );
	OR2X1 U27 ( .A(bouta_fifomodule31), .B(boutb_fifomodule31), .Y(boutmain_fifomodule31) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule31[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule31[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule31) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule31) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(write_ptr_ff_fifomodule31[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(read_ptr_ff_fifomodule31[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(fifo_ff_fifomodule31[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(write_ptr_ff_fifomodule31[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(read_ptr_ff_fifomodule31[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(fifo_ff_fifomodule31[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule31[0]), .Q(write_ptr_ff_fifomodule31[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule31[1]), .Q(write_ptr_ff_fifomodule31[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule31[0]), .Q(read_ptr_ff_fifomodule31[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule31[1]), .Q(read_ptr_ff_fifomodule31[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][0]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][1]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][2]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][3]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][4]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][5]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][6]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][7]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer31), .Y(next_locked_vc_buffer31) );
    BUFX1 U0(.A(flit31[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][0]));
	BUFX1 U1(.A(flit31[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][1]));
	BUFX1 U2(.A(flit31[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][2]));
	BUFX1 U3(.A(flit31[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][3]));
	BUFX1 U4(.A(flit31[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][4]));
	BUFX1 U5(.A(flit31[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][5]));
	BUFX1 U6(.A(flit31[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][6]));
	BUFX1 U7(.A(flit31[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][7]));
	BUFX1 U8(.A(flit31[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][8]));
	BUFX1 U9(.A(flit31[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][9]));
	BUFX1 U10(.A(flit31[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][10]));
	BUFX1 U11(.A(flit31[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][11]));
	BUFX1 U12(.A(flit31[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][12]));
	BUFX1 U13(.A(flit31[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][13]));
	BUFX1 U14(.A(flit31[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][14]));
	BUFX1 U15(.A(flit31[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][15]));
	BUFX1 U16(.A(flit31[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][16]));
	BUFX1 U17(.A(flit31[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][17]));
	BUFX1 U18(.A(flit31[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][18]));
	BUFX1 U19(.A(flit31[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][19]));
	BUFX1 U20(.A(flit31[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][20]));
	BUFX1 U21(.A(flit31[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][21]));
	BUFX1 U22(.A(flit31[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][22]));
	BUFX1 U23(.A(flit31[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][23]));
	BUFX1 U24(.A(flit31[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][24]));
	BUFX1 U25(.A(flit31[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][25]));
	BUFX1 U26(.A(flit31[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][26]));
	BUFX1 U27(.A(flit31[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][27]));
	BUFX1 U28(.A(flit31[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][28]));
	BUFX1 U29(.A(flit31[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][29]));
	BUFX1 U30(.A(flit31[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][30]));
	BUFX1 U31(.A(flit31[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][31]));
	BUFX1 U32(.A(flit31[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][32]));
	BUFX1 U33(.A(flit31[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][33]));
    NOR2X1 U34 ( .IN1(flit31[33]), .IN2(flit31[32]), .QN(norres_vc_buffer31_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit31[29]), .IN2(flit31[28]), .IN3(flit31[27]), .IN4(flit31[26]), .Y(or1res_vc_buffer31) );
    OR4X1 U35 ( .IN1(flit31[25]), .IN2(flit31[24]), .IN3(flit31[23]), .IN4(flit31[22]), .Y(or2res_vc_buffer31) );
    OR2X1 U36 ( .A(or1res_vc_buffer31), .B(or2res_vc_buffer31), .Y(orres_vc_buffer31) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(norres_vc_buffer31_vc_buffer1), .IN3(orres_vc_buffer31), .Q(finres1_vc_buffer31) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer31), .IN2(1'b1), .S(finres1_vc_buffer31), .Q(next_locked_vc_buffer31);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(flit31[33]), .IN3(flit31[32]), .Q(andres1_vc_buffer31) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer31), .IN2(1'b0), .S(andres1_vc_buffer31), .Q(next_locked_vc_buffer31);

    INVX1 U41 ( .A(full_vc_buffer31), .Y(full_vc_buffer31_not1) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer31), .Y(locked_by_route_ff_vc_buffer31_not1) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer31_not1), .S(norres_vc_buffer31_vc_buffer1), .Q(thirdand_vc_buffer31);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(full_vc_buffer31_not1), .IN3(thirdand_vc_buffer31), .Q(write_flit31_vc_buffer13) );
    AND2X1 U45 ( .IN1(full_vc_buffer31_not1), .IN2(norres_vc_buffer31_vc_buffer1), .Q(from_input_resp_input_datapath3[1]) );
    INVX1 U46 ( .A(empty_vc_buffer31), .Y(to_output_req_in_jump_input_datapath3put_datapath3[37]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[37]), .IN2(to_output_resp_input_datapath3[1]), .Q(read_flit31_vc_buffer13) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath3put_datapath3[39:38]), .Y(2'b01));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer31), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer31);


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule32[0]), .Y(next_read_ptr_fifomodule32[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule32[1]), .Y(next_read_ptr_fifomodule32[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule32[0]), .Y(next_write_ptr_fifomodule32[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule32[1]), .Y(next_write_ptr_fifomodule32[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule32[0]), .IN2(read_ptr_ff_fifomodule32[0]), .Q(u1temp_fifomodule32) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule32[1]), .IN2(read_ptr_ff_fifomodule32[1]), .Q(u2temp_fifomodule32) );
	AND2X1 U3 ( .A(u1temp_fifomodule32), .B(u2temp_fifomodule32), .Y(empty_vc_buffer32) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule32[1]), .B(read_ptr_ff_fifomodule32[1]), .Y(u4temp_fifomodule32) );
	AND2X1 U5 ( .A(u1temp_fifomodule32), .B(u4temp_fifomodule32), .Y(full_vc_buffer32) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][7]));

	INVX1 U7 ( .A(full_vc_buffer32), .Y(full_vc_buffer32_not2_fifomodule2) );
	AND2X1 U8 ( .A(write_flit32_vc_buffer23), .B(full_vc_buffer32_not2_fifomodule2), .Y(u7temp_fifomodule32) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule32), .Q(u9temp_fifomodule32));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule32[0]), .B0(u9temp_fifomodule32), .C1(u10carry_fifomodule32), .SO(next_write_ptr_fifomodule32[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule32), .B0(write_ptr_ff_fifomodule32[1]), .C1(u11carry_fifomodule32), .SO(next_write_ptr_fifomodule32[1]) );

	INVX1 U12 ( .A(empty_vc_buffer32), .Y(empty_vc_buffer32_not_fifomodule2) );
	AND2X1 U13 ( .A(read_flit32_vc_buffer23), .B(empty_vc_buffer32_not_fifomodule2), .Y(u13temp_fifomodule32) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule32), .Q(u14temp_fifomodule32));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule32[0]), .B0(u14temp_fifomodule32), .C1(u15carry_fifomodule32), .SO(next_read_ptr_fifomodule32[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule32), .B0(read_ptr_ff_fifomodule32[1]), .C1(u16carry_fifomodule32), .SO(next_read_ptr_fifomodule32[1]) );

	AND2X1 U17 ( .A(write_flit32_vc_buffer23), .B(full_vc_buffer32), .Y(u17res_fifomodule32) );
	AND2X1 U18 ( .A(read_flit32_vc_buffer23), .B(empty_vc_buffer32), .Y(u18res_fifomodule32) );
    OR2X1 U19 ( .A(u17res_fifomodule32), .B(u18res_fifomodule32), .Y(error_vc_buffer32) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule32[0]), .B(read_ptr_ff_fifomodule32[0]), .Y(fifo_ocup_fifomodule32[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule32[0]), .Y(write_ptr_ff_fifomodule32_0_not23) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule32_0_not23), .B(read_ptr_ff_fifomodule32[0]), .Y(b0wire_fifomodule32) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule32[1]), .B(read_ptr_ff_fifomodule32[1]), .Y(u23temp_fifomodule32) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule32[1]), .Y(write_ptr_ff_fifomodule32_1_not23) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule32[1]), .B(write_ptr_ff_fifomodule32_1_not23), .Y(boutb_fifomodule32) );
	XOR2X1 U24 ( .A(u23temp_fifomodule32), .B(b0wire_fifomodule32), .Y(fifo_ocup_fifomodule32[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule32), .Y(u23temp_fifomodule32_not_fifomodule2) );
	AND2X1 U26 ( .A(b0wire_fifomodule32), .B(u23temp_fifomodule32_not_fifomodule2), .Y(bouta_fifomodule32) );
	OR2X1 U27 ( .A(bouta_fifomodule32), .B(boutb_fifomodule32), .Y(boutmain_fifomodule32) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule32[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule32[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule32) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule32) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(write_ptr_ff_fifomodule32[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(read_ptr_ff_fifomodule32[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(fifo_ff_fifomodule32[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(write_ptr_ff_fifomodule32[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(read_ptr_ff_fifomodule32[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(fifo_ff_fifomodule32[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule32[0]), .Q(write_ptr_ff_fifomodule32[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule32[1]), .Q(write_ptr_ff_fifomodule32[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule32[0]), .Q(read_ptr_ff_fifomodule32[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule32[1]), .Q(read_ptr_ff_fifomodule32[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][0]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][1]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][2]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][3]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][4]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][5]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][6]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][7]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer32), .Y(next_locked_vc_buffer32) );
    BUFX1 U0(.A(flit32[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][0]));
	BUFX1 U1(.A(flit32[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][1]));
	BUFX1 U2(.A(flit32[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][2]));
	BUFX1 U3(.A(flit32[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][3]));
	BUFX1 U4(.A(flit32[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][4]));
	BUFX1 U5(.A(flit32[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][5]));
	BUFX1 U6(.A(flit32[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][6]));
	BUFX1 U7(.A(flit32[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][7]));
	BUFX1 U8(.A(flit32[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][8]));
	BUFX1 U9(.A(flit32[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][9]));
	BUFX1 U10(.A(flit32[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][10]));
	BUFX1 U11(.A(flit32[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][11]));
	BUFX1 U12(.A(flit32[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][12]));
	BUFX1 U13(.A(flit32[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][13]));
	BUFX1 U14(.A(flit32[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][14]));
	BUFX1 U15(.A(flit32[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][15]));
	BUFX1 U16(.A(flit32[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][16]));
	BUFX1 U17(.A(flit32[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][17]));
	BUFX1 U18(.A(flit32[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][18]));
	BUFX1 U19(.A(flit32[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][19]));
	BUFX1 U20(.A(flit32[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][20]));
	BUFX1 U21(.A(flit32[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][21]));
	BUFX1 U22(.A(flit32[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][22]));
	BUFX1 U23(.A(flit32[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][23]));
	BUFX1 U24(.A(flit32[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][24]));
	BUFX1 U25(.A(flit32[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][25]));
	BUFX1 U26(.A(flit32[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][26]));
	BUFX1 U27(.A(flit32[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][27]));
	BUFX1 U28(.A(flit32[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][28]));
	BUFX1 U29(.A(flit32[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][29]));
	BUFX1 U30(.A(flit32[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][30]));
	BUFX1 U31(.A(flit32[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][31]));
	BUFX1 U32(.A(flit32[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][32]));
	BUFX1 U33(.A(flit32[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][33]));
    NOR2X1 U34 ( .IN1(flit32[33]), .IN2(flit32[32]), .QN(norres_vc_buffer32_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit32[29]), .IN2(flit32[28]), .IN3(flit32[27]), .IN4(flit32[26]), .Y(or1res_vc_buffer32) );
    OR4X1 U35 ( .IN1(flit32[25]), .IN2(flit32[24]), .IN3(flit32[23]), .IN4(flit32[22]), .Y(or2res_vc_buffer32) );
    OR2X1 U36 ( .A(or1res_vc_buffer32), .B(or2res_vc_buffer32), .Y(orres_vc_buffer32) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(norres_vc_buffer32_vc_buffer2), .IN3(orres_vc_buffer32), .Q(finres1_vc_buffer32) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer32), .IN2(1'b1), .S(finres1_vc_buffer32), .Q(next_locked_vc_buffer32);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(flit32[33]), .IN3(flit32[32]), .Q(andres1_vc_buffer32) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer32), .IN2(1'b0), .S(andres1_vc_buffer32), .Q(next_locked_vc_buffer32);

    INVX1 U41 ( .A(full_vc_buffer32), .Y(full_vc_buffer32_not2) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer32), .Y(locked_by_route_ff_vc_buffer32_not2) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer32_not2), .S(norres_vc_buffer32_vc_buffer2), .Q(thirdand_vc_buffer32);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(full_vc_buffer32_not2), .IN3(thirdand_vc_buffer32), .Q(write_flit32_vc_buffer23) );
    AND2X1 U45 ( .IN1(full_vc_buffer32_not2), .IN2(norres_vc_buffer32_vc_buffer2), .Q(from_input_resp_input_datapath3[2]) );
    INVX1 U46 ( .A(empty_vc_buffer32), .Y(to_output_req_in_jump_input_datapath3put_datapath3[74]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[74]), .IN2(to_output_resp_input_datapath3[2]), .Q(read_flit32_vc_buffer23) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath3put_datapath3[76:75]), .Y(2'b10));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer32), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer32);

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath3put_datapath3[77]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath3put_datapath3[78]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath3put_datapath3[79]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath3put_datapath3[80]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath3put_datapath3[81]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath3put_datapath3[82]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath3put_datapath3[83]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath3put_datapath3[84]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath3put_datapath3[85]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath3put_datapath3[86]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath3put_datapath3[87]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath3put_datapath3[88]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath3put_datapath3[89]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath3put_datapath3[90]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath3put_datapath3[91]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath3put_datapath3[92]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath3put_datapath3[93]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath3put_datapath3[94]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath3put_datapath3[95]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath3put_datapath3[96]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath3put_datapath3[97]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath3put_datapath3[98]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath3put_datapath3[99]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath3put_datapath3[100]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath3put_datapath3[101]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath3put_datapath3[102]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath3put_datapath3[103]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath3put_datapath3[104]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath3put_datapath3[105]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath3put_datapath3[106]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath3put_datapath3[107]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath3put_datapath3[108]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath3put_datapath3[109]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath3put_datapath3[110]), .Y(ext_req_v_i[147:111][36]));
    XNOR2X1 U222 ( .IN1(ext_req_v_i[147:111][1]), .IN2(i_input_datapath3[0]), .QN(xnor1resu_input_datapath3) );
    XNOR2X1 U222 ( .IN1(ext_req_v_i[147:111][2]), .IN2(i_input_datapath3[1]), .QN(xnor2resu_input_datapath3) );
    AND2X1 U128 ( .IN1(xnor1resu_input_datapath3), .IN2(xnor2resu_input_datapath3), .Q(and1resu_input_datapath3) );
    AND3X1 U128 ( .IN1(and1resu_input_datapath3), .IN2(ext_req_v_i[147:111][0]), .IN2(ext_req_v_i[147:111][0]), .Q(cond1line_input_datapath3) );
    MUX21X1 U0009 (.IN1(vc_ch_act_in_input_datapath3[0]), .IN2(i_input_datapath3[0]), .S(cond1line_input_datapath3), .Q(vc_ch_act_in_input_datapath3[0]));
    MUX21X1 U0010 (.IN1(vc_ch_act_in_input_datapath3[1]), .IN2(i_input_datapath3[1]), .S(cond1line_input_datapath3), .Q(vc_ch_act_in_input_datapath3[1]));
    MUX21X1 U0011 (.IN1(req_in_jump_input_datapath3), .IN2(1), .S(cond1line_input_datapath3), .Q(req_in_jump_input_datapath3));
	BUFX1 U3(.A(from_input_req_in_jump_input_datapath3put_datapath3[40]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath3put_datapath3[41]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath3put_datapath3[42]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath3put_datapath3[43]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath3put_datapath3[44]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath3put_datapath3[45]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath3put_datapath3[46]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath3put_datapath3[47]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath3put_datapath3[48]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath3put_datapath3[49]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath3put_datapath3[50]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath3put_datapath3[51]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath3put_datapath3[52]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath3put_datapath3[53]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath3put_datapath3[54]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath3put_datapath3[55]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath3put_datapath3[56]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath3put_datapath3[57]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath3put_datapath3[58]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath3put_datapath3[59]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath3put_datapath3[60]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath3put_datapath3[61]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath3put_datapath3[62]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath3put_datapath3[63]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath3put_datapath3[64]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath3put_datapath3[65]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath3put_datapath3[66]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath3put_datapath3[67]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath3put_datapath3[68]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath3put_datapath3[69]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath3put_datapath3[70]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath3put_datapath3[71]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath3put_datapath3[72]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath3put_datapath3[73]), .Y(ext_req_v_i[147:111][36]));

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath3put_datapath3[3]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath3put_datapath3[4]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath3put_datapath3[5]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath3put_datapath3[6]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath3put_datapath3[7]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath3put_datapath3[8]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath3put_datapath3[9]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath3put_datapath3[10]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath3put_datapath3[11]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath3put_datapath3[12]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath3put_datapath3[13]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath3put_datapath3[14]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath3put_datapath3[15]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath3put_datapath3[16]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath3put_datapath3[17]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath3put_datapath3[18]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath3put_datapath3[19]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath3put_datapath3[20]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath3put_datapath3[21]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath3put_datapath3[22]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath3put_datapath3[23]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath3put_datapath3[24]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath3put_datapath3[25]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath3put_datapath3[26]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath3put_datapath3[27]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath3put_datapath3[28]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath3put_datapath3[29]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath3put_datapath3[30]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath3put_datapath3[31]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath3put_datapath3[32]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath3put_datapath3[33]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath3put_datapath3[34]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath3put_datapath3[35]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath3put_datapath3[36]), .Y(ext_req_v_i[147:111][36]));

    MUX21X1 U0012 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3 * 37]), .IN2(ext_req_v_i[147:111][0]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3 * 37]));
    MUX21X1 U0013 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+2]), .IN2(vc_ch_act_in_input_datapath3[1]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+2]));
    MUX21X1 U0014 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+1]), .IN2(vc_ch_act_in_input_datapath3[0]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+1]));
    MUX21X1 U0015 (.IN1(ext_resp_v_o[4:3][0]), .IN2(from_input_resp_input_datapath3[vc_ch_act_in_input_datapath3]), .S(req_in_jump_input_datapath3), .Q(ext_resp_v_o[4:3][0]));

    INVX1 U041 ( .A(req_in_jump_input_datapath3), .Y(req_in_jump_input_datapath3_not) );
    MUX21X1 U0016 (.IN1(ext_resp_v_o[4:3][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath3_not), .Q(ext_resp_v_o[4:3][0]));
    BUFX1 U34(.A(from_input_req_in_jump_input_datapath3put_datapath3[34]), .Y(ext_req_v_i[147:111][34]));

    XOR2X1 U0222 ( .IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b1), .Q(xor1resu_input_datapath3) );
    MUX21X1 U0017 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(xor1resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U0018 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b0), .S(xor1resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[1]));
    AND2X1 U38123 ( .IN1(xor1resu_input_datapath3), .IN2(to_output_req_in_jump_input_datapath3put_datapath3[j_input_datapath3*37]), .Q(and2resu_input_datapath3) );
    MUX21X1 U0019 (.IN1(vc_ch_act_out_input_datapath3[0]), .IN2(j_input_datapath3[0]), .S(and2resu_input_datapath3), .Q(vc_ch_act_out_input_datapath3[0]));
    MUX21X1 U0020 (.IN1(vc_ch_act_out_input_datapath3[1]), .IN2(j_input_datapath3[1]), .S(and2resu_input_datapath3), .Q(vc_ch_act_out_input_datapath3[1]));
    MUX21X1 U0021 (.IN1(req_out_jump_input_datapath3), .IN2(1'b1), .S(and2resu_input_datapath3), .Q(req_out_jump_input_datapath3));
    MUX21X1 U0022 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(and2resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U0023 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b1), .S(and2resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[1]));
    HADDX1 U00021 ( .A0(j_input_datapath3[0]), .B0(1'b1), .C1(j_input_datapath3[1]), .SO(j_input_datapath3[0]) );
    HADDX1 U00022 ( .A0(j_input_datapath3[0]), .B0(1'b1), .C1(j_input_datapath3[1]), .SO(j_input_datapath3[0]) );
    AND2X1 U38111 ( .IN1(xor1resu_input_datapath3), .IN2(to_output_req_in_jump_input_datapath3put_datapath3[j_input_datapath3*37]), .Q(and3resu) );
    NAND2X1 U29311(.A(_sv2v_jump_input_datapath3[0]),.B(_sv2v_jump_input_datapath3[1]),.Y(nand1resu_input_datapath33));
    MUX21X1 U00212 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(nand1resu_input_datapath33), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U00213 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b0), .S(nand1resu_input_datapath33), .Q(_sv2v_jump_input_datapath3[1]));
    XNOR2X1 U17581 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(_sv2v_jump_input_datapath3[1]), .Q(xnor23resu_input_datapath3) );
    AND2X1 U38111 ( .IN1(xnor23resu_input_datapath3), .IN2(req_out_jump_input_datapath3), .Q(and4resu_input_datapath3) );

    MUX21X1 U3(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[147:111][3]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U4(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[147:111][4]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U5(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[147:111][5]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U6(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[147:111][6]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U7(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[147:111][7]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U8(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[147:111][8]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U9(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[147:111][9]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U10(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[147:111][10]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U11(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[147:111][11]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U12(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[147:111][12]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U13(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[147:111][13]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U14(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[147:111][14]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U15(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[147:111][15]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U16(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[147:111][16]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U17(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[147:111][17]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U18(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[147:111][18]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U19(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[147:111][19]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U20(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[147:111][20]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U21(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[147:111][21]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U22(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[147:111][22]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U23(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[147:111][23]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U24(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[147:111][24]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U25(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[147:111][25]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U26(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[147:111][26]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U27(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[147:111][27]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U28(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[147:111][28]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U29(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[147:111][29]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U30(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[147:111][30]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U31(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[147:111][31]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U32(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[147:111][32]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U33(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[147:111][33]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U34(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[147:111][34]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U35(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[147:111][35]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U36(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[147:111][36]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U321111(.IN1(int_req_v[147:111][0]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3 * 37)]), .S(and4resu_input_datapath3), .Q(int_req_v[147:111][0]));
	MUX21X1 U331112(.IN1(int_req_v[147:111][1]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+1]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+1]));
	MUX21X1 U331122(.IN1(int_req_v[147:111][2]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+2]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3]),.IN2(int_resp_v[4:3]), .S(and4resu_input_datapath3), .Q(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3+1]),.IN2(int_resp_v[4:3]), .S(and4resu_input_datapath3), .Q(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3+1]));

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule4[0]), .Y(next_read_ptr_fifomodule4[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule4[1]), .Y(next_read_ptr_fifomodule4[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule4[0]), .Y(next_write_ptr_fifomodule4[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule4[1]), .Y(next_write_ptr_fifomodule4[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule4[0]), .IN2(read_ptr_ff_fifomodule4[0]), .Q(u1temp_fifomodule4) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule4[1]), .IN2(read_ptr_ff_fifomodule4[1]), .Q(u2temp_fifomodule4) );
	AND2X1 U3 ( .A(u1temp_fifomodule4), .B(u2temp_fifomodule4), .Y(empty_vc_buffer4) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule4[1]), .B(read_ptr_ff_fifomodule4[1]), .Y(u4temp_fifomodule4) );
	AND2X1 U5 ( .A(u1temp_fifomodule4), .B(u4temp_fifomodule4), .Y(full_vc_buffer4) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][7]));

	INVX1 U7 ( .A(full_vc_buffer4), .Y(full_vc_buffer4_not_fifomodule) );
	AND2X1 U8 ( .A(write_flit4_vc_buffer4), .B(full_vc_buffer4_not_fifomodule), .Y(u7temp_fifomodule4) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule4), .Q(u9temp_fifomodule4));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule4[0]), .B0(u9temp_fifomodule4), .C1(u10carry_fifomodule4), .SO(next_write_ptr_fifomodule4[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule4), .B0(write_ptr_ff_fifomodule4[1]), .C1(u11carry_fifomodule4), .SO(next_write_ptr_fifomodule4[1]) );

	INVX1 U12 ( .A(empty_vc_buffer4), .Y(empty_vc_buffer4_not_fifomodule) );
	AND2X1 U13 ( .A(read_flit4_vc_buffer4), .B(empty_vc_buffer4_not_fifomodule), .Y(u13temp_fifomodule4) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule4), .Q(u14temp_fifomodule4));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule4[0]), .B0(u14temp_fifomodule4), .C1(u15carry_fifomodule4), .SO(next_read_ptr_fifomodule4[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule4), .B0(read_ptr_ff_fifomodule4[1]), .C1(u16carry_fifomodule4), .SO(next_read_ptr_fifomodule4[1]) );

	AND2X1 U17 ( .A(write_flit4_vc_buffer4), .B(full_vc_buffer4), .Y(u17res_fifomodule4) );
	AND2X1 U18 ( .A(read_flit4_vc_buffer4), .B(empty_vc_buffer4), .Y(u18res_fifomodule4) );
    OR2X1 U19 ( .A(u17res_fifomodule4), .B(u18res_fifomodule4), .Y(error_vc_buffer4) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule4[0]), .B(read_ptr_ff_fifomodule4[0]), .Y(fifo_ocup_fifomodule4[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule4[0]), .Y(write_ptr_ff_fifomodule4_0_not4) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule4_0_not4), .B(read_ptr_ff_fifomodule4[0]), .Y(b0wire_fifomodule4) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule4[1]), .B(read_ptr_ff_fifomodule4[1]), .Y(u23temp_fifomodule4) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule4[1]), .Y(write_ptr_ff_fifomodule4_1_not4) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule4[1]), .B(write_ptr_ff_fifomodule4_1_not4), .Y(boutb_fifomodule4) );
	XOR2X1 U24 ( .A(u23temp_fifomodule4), .B(b0wire_fifomodule4), .Y(fifo_ocup_fifomodule4[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule4), .Y(u23temp_fifomodule4_not_fifomodule4) );
	AND2X1 U26 ( .A(b0wire_fifomodule4), .B(u23temp_fifomodule4_not_fifomodule4), .Y(bouta_fifomodule4) );
	OR2X1 U27 ( .A(bouta_fifomodule4), .B(boutb_fifomodule4), .Y(boutmain_fifomodule4) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule4[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule4[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule4) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule4) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(write_ptr_ff_fifomodule4[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(read_ptr_ff_fifomodule4[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(fifo_ff_fifomodule4[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(write_ptr_ff_fifomodule4[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(read_ptr_ff_fifomodule4[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(fifo_ff_fifomodule4[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule4[0]), .Q(write_ptr_ff_fifomodule4[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule4[1]), .Q(write_ptr_ff_fifomodule4[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule4[0]), .Q(read_ptr_ff_fifomodule4[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule4[1]), .Q(read_ptr_ff_fifomodule4[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][0]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][1]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][2]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][3]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][4]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][5]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][6]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][7]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer4), .Y(next_locked_vc_buffer4) );
    BUFX1 U0(.A(flit4[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][0]));
	BUFX1 U1(.A(flit4[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][1]));
	BUFX1 U2(.A(flit4[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][2]));
	BUFX1 U3(.A(flit4[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][3]));
	BUFX1 U4(.A(flit4[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][4]));
	BUFX1 U5(.A(flit4[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][5]));
	BUFX1 U6(.A(flit4[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][6]));
	BUFX1 U7(.A(flit4[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][7]));
	BUFX1 U8(.A(flit4[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][8]));
	BUFX1 U9(.A(flit4[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][9]));
	BUFX1 U10(.A(flit4[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][10]));
	BUFX1 U11(.A(flit4[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][11]));
	BUFX1 U12(.A(flit4[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][12]));
	BUFX1 U13(.A(flit4[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][13]));
	BUFX1 U14(.A(flit4[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][14]));
	BUFX1 U15(.A(flit4[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][15]));
	BUFX1 U16(.A(flit4[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][16]));
	BUFX1 U17(.A(flit4[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][17]));
	BUFX1 U18(.A(flit4[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][18]));
	BUFX1 U19(.A(flit4[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][19]));
	BUFX1 U20(.A(flit4[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][20]));
	BUFX1 U21(.A(flit4[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][21]));
	BUFX1 U22(.A(flit4[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][22]));
	BUFX1 U23(.A(flit4[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][23]));
	BUFX1 U24(.A(flit4[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][24]));
	BUFX1 U25(.A(flit4[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][25]));
	BUFX1 U26(.A(flit4[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][26]));
	BUFX1 U27(.A(flit4[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][27]));
	BUFX1 U28(.A(flit4[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][28]));
	BUFX1 U29(.A(flit4[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][29]));
	BUFX1 U30(.A(flit4[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][30]));
	BUFX1 U31(.A(flit4[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][31]));
	BUFX1 U32(.A(flit4[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][32]));
	BUFX1 U33(.A(flit4[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][33]));
    NOR2X1 U34 ( .IN1(flit4[33]), .IN2(flit4[32]), .QN(norres_vc_buffer4_vc_buffer4) );
    OR4X1 U35 ( .IN1(flit4[29]), .IN2(flit4[28]), .IN3(flit4[27]), .IN4(flit4[26]), .Y(or1res_vc_buffer4) );
    OR4X1 U35 ( .IN1(flit4[25]), .IN2(flit4[24]), .IN3(flit4[23]), .IN4(flit4[22]), .Y(or2res_vc_buffer4) );
    OR2X1 U36 ( .A(or1res_vc_buffer4), .B(or2res_vc_buffer4), .Y(orres_vc_buffer4) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(norres_vc_buffer4_vc_buffer4), .IN3(orres_vc_buffer4), .Q(finres1_vc_buffer4) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer4), .IN2(1'b1), .S(finres1_vc_buffer4), .Q(next_locked_vc_buffer4);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(flit4[33]), .IN3(flit4[32]), .Q(andres1_vc_buffer4) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer4), .IN2(1'b0), .S(andres1_vc_buffer4), .Q(next_locked_vc_buffer4);

    INVX1 U41 ( .A(full_vc_buffer4), .Y(full_vc_buffer4_not) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer4), .Y(locked_by_route_ff_vc_buffer4_not) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer4_not), .S(norres_vc_buffer4_vc_buffer4), .Q(thirdand_vc_buffer4);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(full_vc_buffer4_not), .IN3(thirdand_vc_buffer4), .Q(write_flit4_vc_buffer4) );
    AND2X1 U45 ( .IN1(full_vc_buffer4_not), .IN2(norres_vc_buffer4_vc_buffer4), .Q(from_input_resp_input_datapath4[0]) );
    INVX1 U46 ( .A(empty_vc_buffer4), .Y(to_output_req_in_jump_input_datapath4put_datapath4[0]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[0]), .IN2(to_output_resp_input_datapath4[0]), .Q(read_flit4_vc_buffer4) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath4put_datapath4[2:1]), .Y(2'b00));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer4), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer4);

	BUFX1 U00 ( .A(read_ptr_ff_fifomodule41[0]), .Y(next_read_ptr_fifomodule41[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule41[1]), .Y(next_read_ptr_fifomodule41[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule41[0]), .Y(next_write_ptr_fifomodule41[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule41[1]), .Y(next_write_ptr_fifomodule41[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule41[0]), .IN2(read_ptr_ff_fifomodule41[0]), .Q(u1temp_fifomodule41) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule41[1]), .IN2(read_ptr_ff_fifomodule41[1]), .Q(u2temp_fifomodule41) );
	AND2X1 U3 ( .A(u1temp_fifomodule41), .B(u2temp_fifomodule41), .Y(empty_vc_buffer41) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule41[1]), .B(read_ptr_ff_fifomodule41[1]), .Y(u4temp_fifomodule41) );
	AND2X1 U5 ( .A(u1temp_fifomodule41), .B(u4temp_fifomodule41), .Y(full_vc_buffer41) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][7]));

	INVX1 U7 ( .A(full_vc_buffer41), .Y(full_vc_buffer41_not1_fifomodule1) );
	AND2X1 U8 ( .A(write_flit41_vc_buffer14), .B(full_vc_buffer41_not1_fifomodule1), .Y(u7temp_fifomodule41) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule41), .Q(u9temp_fifomodule41));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule41[0]), .B0(u9temp_fifomodule41), .C1(u10carry_fifomodule41), .SO(next_write_ptr_fifomodule41[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule41), .B0(write_ptr_ff_fifomodule41[1]), .C1(u11carry_fifomodule41), .SO(next_write_ptr_fifomodule41[1]) );

	INVX1 U12 ( .A(empty_vc_buffer41), .Y(empty_vc_buffer41_not_fifomodule1) );
	AND2X1 U13 ( .A(read_flit41_vc_buffer14), .B(empty_vc_buffer41_not_fifomodule1), .Y(u13temp_fifomodule41) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule41), .Q(u14temp_fifomodule41));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule41[0]), .B0(u14temp_fifomodule41), .C1(u15carry_fifomodule41), .SO(next_read_ptr_fifomodule41[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule41), .B0(read_ptr_ff_fifomodule41[1]), .C1(u16carry_fifomodule41), .SO(next_read_ptr_fifomodule41[1]) );

	AND2X1 U17 ( .A(write_flit41_vc_buffer14), .B(full_vc_buffer41), .Y(u17res_fifomodule41) );
	AND2X1 U18 ( .A(read_flit41_vc_buffer14), .B(empty_vc_buffer41), .Y(u18res_fifomodule41) );
    OR2X1 U19 ( .A(u17res_fifomodule41), .B(u18res_fifomodule41), .Y(error_vc_buffer41) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule41[0]), .B(read_ptr_ff_fifomodule41[0]), .Y(fifo_ocup_fifomodule41[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule41[0]), .Y(write_ptr_ff_fifomodule41_0_not14) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule41_0_not14), .B(read_ptr_ff_fifomodule41[0]), .Y(b0wire_fifomodule41) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule41[1]), .B(read_ptr_ff_fifomodule41[1]), .Y(u23temp_fifomodule41) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule41[1]), .Y(write_ptr_ff_fifomodule41_1_not14) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule41[1]), .B(write_ptr_ff_fifomodule41_1_not14), .Y(boutb_fifomodule41) );
	XOR2X1 U24 ( .A(u23temp_fifomodule41), .B(b0wire_fifomodule41), .Y(fifo_ocup_fifomodule41[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule41), .Y(u23temp_fifomodule41_not_fifomodule1) );
	AND2X1 U26 ( .A(b0wire_fifomodule41), .B(u23temp_fifomodule41_not_fifomodule1), .Y(bouta_fifomodule41) );
	OR2X1 U27 ( .A(bouta_fifomodule41), .B(boutb_fifomodule41), .Y(boutmain_fifomodule41) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule41[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule41[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule41) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule41) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(write_ptr_ff_fifomodule41[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(read_ptr_ff_fifomodule41[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(fifo_ff_fifomodule41[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(write_ptr_ff_fifomodule41[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(read_ptr_ff_fifomodule41[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(fifo_ff_fifomodule41[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule41[0]), .Q(write_ptr_ff_fifomodule41[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule41[1]), .Q(write_ptr_ff_fifomodule41[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule41[0]), .Q(read_ptr_ff_fifomodule41[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule41[1]), .Q(read_ptr_ff_fifomodule41[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][0]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][1]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][2]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][3]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][4]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][5]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][6]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][7]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer41), .Y(next_locked_vc_buffer41) );
    BUFX1 U0(.A(flit41[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][0]));
	BUFX1 U1(.A(flit41[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][1]));
	BUFX1 U2(.A(flit41[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][2]));
	BUFX1 U3(.A(flit41[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][3]));
	BUFX1 U4(.A(flit41[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][4]));
	BUFX1 U5(.A(flit41[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][5]));
	BUFX1 U6(.A(flit41[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][6]));
	BUFX1 U7(.A(flit41[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][7]));
	BUFX1 U8(.A(flit41[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][8]));
	BUFX1 U9(.A(flit41[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][9]));
	BUFX1 U10(.A(flit41[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][10]));
	BUFX1 U11(.A(flit41[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][11]));
	BUFX1 U12(.A(flit41[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][12]));
	BUFX1 U13(.A(flit41[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][13]));
	BUFX1 U14(.A(flit41[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][14]));
	BUFX1 U15(.A(flit41[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][15]));
	BUFX1 U16(.A(flit41[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][16]));
	BUFX1 U17(.A(flit41[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][17]));
	BUFX1 U18(.A(flit41[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][18]));
	BUFX1 U19(.A(flit41[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][19]));
	BUFX1 U20(.A(flit41[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][20]));
	BUFX1 U21(.A(flit41[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][21]));
	BUFX1 U22(.A(flit41[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][22]));
	BUFX1 U23(.A(flit41[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][23]));
	BUFX1 U24(.A(flit41[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][24]));
	BUFX1 U25(.A(flit41[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][25]));
	BUFX1 U26(.A(flit41[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][26]));
	BUFX1 U27(.A(flit41[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][27]));
	BUFX1 U28(.A(flit41[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][28]));
	BUFX1 U29(.A(flit41[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][29]));
	BUFX1 U30(.A(flit41[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][30]));
	BUFX1 U31(.A(flit41[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][31]));
	BUFX1 U32(.A(flit41[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][32]));
	BUFX1 U33(.A(flit41[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][33]));
    NOR2X1 U34 ( .IN1(flit41[33]), .IN2(flit41[32]), .QN(norres_vc_buffer41_vc_buffer1) );
    OR4X1 U35 ( .IN1(flit41[29]), .IN2(flit41[28]), .IN3(flit41[27]), .IN4(flit41[26]), .Y(or1res_vc_buffer41) );
    OR4X1 U35 ( .IN1(flit41[25]), .IN2(flit41[24]), .IN3(flit41[23]), .IN4(flit41[22]), .Y(or2res_vc_buffer41) );
    OR2X1 U36 ( .A(or1res_vc_buffer41), .B(or2res_vc_buffer41), .Y(orres_vc_buffer41) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(norres_vc_buffer41_vc_buffer1), .IN3(orres_vc_buffer41), .Q(finres1_vc_buffer41) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer41), .IN2(1'b1), .S(finres1_vc_buffer41), .Q(next_locked_vc_buffer41);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(flit41[33]), .IN3(flit41[32]), .Q(andres1_vc_buffer41) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer41), .IN2(1'b0), .S(andres1_vc_buffer41), .Q(next_locked_vc_buffer41);

    INVX1 U41 ( .A(full_vc_buffer41), .Y(full_vc_buffer41_not1) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer41), .Y(locked_by_route_ff_vc_buffer41_not1) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer41_not1), .S(norres_vc_buffer41_vc_buffer1), .Q(thirdand_vc_buffer41);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(full_vc_buffer41_not1), .IN3(thirdand_vc_buffer41), .Q(write_flit41_vc_buffer14) );
    AND2X1 U45 ( .IN1(full_vc_buffer41_not1), .IN2(norres_vc_buffer41_vc_buffer1), .Q(from_input_resp_input_datapath4[1]) );
    INVX1 U46 ( .A(empty_vc_buffer41), .Y(to_output_req_in_jump_input_datapath4put_datapath4[37]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[37]), .IN2(to_output_resp_input_datapath4[1]), .Q(read_flit41_vc_buffer14) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath4put_datapath4[39:38]), .Y(2'b01));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer41), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer41);


	BUFX1 U00 ( .A(read_ptr_ff_fifomodule42[0]), .Y(next_read_ptr_fifomodule42[0]) );
	BUFX1 U01 ( .A(read_ptr_ff_fifomodule42[1]), .Y(next_read_ptr_fifomodule42[1]) );
	BUFX1 U02 ( .A(write_ptr_ff_fifomodule42[0]), .Y(next_write_ptr_fifomodule42[0]) );
	BUFX1 U03 ( .A(write_ptr_ff_fifomodule42[1]), .Y(next_write_ptr_fifomodule42[1]) );

	XNOR2X1 U1 ( .IN1(write_ptr_ff_fifomodule42[0]), .IN2(read_ptr_ff_fifomodule42[0]), .Q(u1temp_fifomodule42) );
	XNOR2X1 U2 ( .IN1(write_ptr_ff_fifomodule42[1]), .IN2(read_ptr_ff_fifomodule42[1]), .Q(u2temp_fifomodule42) );
	AND2X1 U3 ( .A(u1temp_fifomodule42), .B(u2temp_fifomodule42), .Y(empty_vc_buffer42) );
	XOR2X1 U4 ( .A(write_ptr_ff_fifomodule42[1]), .B(read_ptr_ff_fifomodule42[1]), .Y(u4temp_fifomodule42) );
	AND2X1 U5 ( .A(u1temp_fifomodule42), .B(u4temp_fifomodule42), .Y(full_vc_buffer42) );
	MUX21X1 U6 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][0]));
	MUX21X1 U61 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][1]));
	MUX21X1 U62 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][2]));
	MUX21X1 U63 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][3]));
	MUX21X1 U64 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][4]));
	MUX21X1 U65 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][5]));
	MUX21X1 U66 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][6]));
	MUX21X1 U67 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][7]));

	INVX1 U7 ( .A(full_vc_buffer42), .Y(full_vc_buffer42_not2_fifomodule2) );
	AND2X1 U8 ( .A(write_flit42_vc_buffer24), .B(full_vc_buffer42_not2_fifomodule2), .Y(u7temp_fifomodule42) );
	MUX21X1 U9 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule42), .Q(u9temp_fifomodule42));
	HADDX1 U10 ( .A0(write_ptr_ff_fifomodule42[0]), .B0(u9temp_fifomodule42), .C1(u10carry_fifomodule42), .SO(next_write_ptr_fifomodule42[0]) );
	HADDX1 U11 ( .A0(u10carry_fifomodule42), .B0(write_ptr_ff_fifomodule42[1]), .C1(u11carry_fifomodule42), .SO(next_write_ptr_fifomodule42[1]) );

	INVX1 U12 ( .A(empty_vc_buffer42), .Y(empty_vc_buffer42_not_fifomodule2) );
	AND2X1 U13 ( .A(read_flit42_vc_buffer24), .B(empty_vc_buffer42_not_fifomodule2), .Y(u13temp_fifomodule42) );
	MUX21X1 U14 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule42), .Q(u14temp_fifomodule42));
	HADDX1 U15 ( .A0(read_ptr_ff_fifomodule42[0]), .B0(u14temp_fifomodule42), .C1(u15carry_fifomodule42), .SO(next_read_ptr_fifomodule42[0]) );
	HADDX1 U16 ( .A0(u15carry_fifomodule42), .B0(read_ptr_ff_fifomodule42[1]), .C1(u16carry_fifomodule42), .SO(next_read_ptr_fifomodule42[1]) );

	AND2X1 U17 ( .A(write_flit42_vc_buffer24), .B(full_vc_buffer42), .Y(u17res_fifomodule42) );
	AND2X1 U18 ( .A(read_flit42_vc_buffer24), .B(empty_vc_buffer42), .Y(u18res_fifomodule42) );
    OR2X1 U19 ( .A(u17res_fifomodule42), .B(u18res_fifomodule42), .Y(error_vc_buffer42) );
	XOR2X1 U20 ( .A(write_ptr_ff_fifomodule42[0]), .B(read_ptr_ff_fifomodule42[0]), .Y(fifo_ocup_fifomodule42[0]) );
	INVX1 U21 ( .A(write_ptr_ff_fifomodule42[0]), .Y(write_ptr_ff_fifomodule42_0_not24) );
	AND2X1 U22 ( .A(write_ptr_ff_fifomodule42_0_not24), .B(read_ptr_ff_fifomodule42[0]), .Y(b0wire_fifomodule42) );
	XOR2X1 U23 ( .A(write_ptr_ff_fifomodule42[1]), .B(read_ptr_ff_fifomodule42[1]), .Y(u23temp_fifomodule42) );
	INVX1 U24 ( .A(write_ptr_ff_fifomodule42[1]), .Y(write_ptr_ff_fifomodule42_1_not24) );
	AND2X1 U25 ( .A(read_ptr_ff_fifomodule42[1]), .B(write_ptr_ff_fifomodule42_1_not24), .Y(boutb_fifomodule42) );
	XOR2X1 U24 ( .A(u23temp_fifomodule42), .B(b0wire_fifomodule42), .Y(fifo_ocup_fifomodule42[1]) );
	INVX1 U25 ( .A(u23temp_fifomodule42), .Y(u23temp_fifomodule42_not_fifomodule2) );
	AND2X1 U26 ( .A(b0wire_fifomodule42), .B(u23temp_fifomodule42_not_fifomodule2), .Y(bouta_fifomodule42) );
	OR2X1 U27 ( .A(bouta_fifomodule42), .B(boutb_fifomodule42), .Y(boutmain_fifomodule42) );
	DFFX2 U28 ( .CLK(clk), .D(fifo_ocup_fifomodule42[0]), .Q(ocup_o[0]) );
	DFFX2 U29 ( .CLK(clk), .D(fifo_ocup_fifomodule42[1]), .Q(ocup_o[1]) );
	DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule42) );
	DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule42) );
	DFFX2 U32 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(write_ptr_ff_fifomodule42[0]) );
	DFFX2 U33 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(read_ptr_ff_fifomodule42[0]) );
	DFFX2 U34 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(fifo_ff_fifomodule42[0]) );
	DFFX2 U35 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(write_ptr_ff_fifomodule42[1]) );
	DFFX2 U36 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(read_ptr_ff_fifomodule42[1]) );
	DFFX2 U37 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(fifo_ff_fifomodule42[1]) );

	DFFX2 U38 ( .CLK(clk), .D(next_write_ptr_fifomodule42[0]), .Q(write_ptr_ff_fifomodule42[0]) );
	DFFX2 U39 ( .CLK(clk), .D(next_write_ptr_fifomodule42[1]), .Q(write_ptr_ff_fifomodule42[1]) );
	DFFX2 U40 ( .CLK(clk), .D(next_read_ptr_fifomodule42[0]), .Q(read_ptr_ff_fifomodule42[0]) );
	DFFX2 U41 ( .CLK(clk), .D(next_read_ptr_fifomodule42[1]), .Q(read_ptr_ff_fifomodule42[1]) );
	  

	DFFX2 U42 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][0]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8]) );
	DFFX2 U43 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][1]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+1]) );
	DFFX2 U44 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][2]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+2]) );
	DFFX2 U45 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][3]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+3]) );
	DFFX2 U46 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][4]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+4]) );
	DFFX2 U47 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][5]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+5]) );
	DFFX2 U48 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][6]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+6]) );
	DFFX2 U49 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][7]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+7]) );

    BUFX1 U00 ( .A(locked_by_route_ff_vc_buffer42), .Y(next_locked_vc_buffer42) );
    BUFX1 U0(.A(flit42[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][0]));
	BUFX1 U1(.A(flit42[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][1]));
	BUFX1 U2(.A(flit42[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][2]));
	BUFX1 U3(.A(flit42[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][3]));
	BUFX1 U4(.A(flit42[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][4]));
	BUFX1 U5(.A(flit42[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][5]));
	BUFX1 U6(.A(flit42[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][6]));
	BUFX1 U7(.A(flit42[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][7]));
	BUFX1 U8(.A(flit42[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][8]));
	BUFX1 U9(.A(flit42[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][9]));
	BUFX1 U10(.A(flit42[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][10]));
	BUFX1 U11(.A(flit42[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][11]));
	BUFX1 U12(.A(flit42[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][12]));
	BUFX1 U13(.A(flit42[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][13]));
	BUFX1 U14(.A(flit42[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][14]));
	BUFX1 U15(.A(flit42[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][15]));
	BUFX1 U16(.A(flit42[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][16]));
	BUFX1 U17(.A(flit42[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][17]));
	BUFX1 U18(.A(flit42[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][18]));
	BUFX1 U19(.A(flit42[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][19]));
	BUFX1 U20(.A(flit42[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][20]));
	BUFX1 U21(.A(flit42[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][21]));
	BUFX1 U22(.A(flit42[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][22]));
	BUFX1 U23(.A(flit42[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][23]));
	BUFX1 U24(.A(flit42[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][24]));
	BUFX1 U25(.A(flit42[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][25]));
	BUFX1 U26(.A(flit42[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][26]));
	BUFX1 U27(.A(flit42[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][27]));
	BUFX1 U28(.A(flit42[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][28]));
	BUFX1 U29(.A(flit42[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][29]));
	BUFX1 U30(.A(flit42[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][30]));
	BUFX1 U31(.A(flit42[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][31]));
	BUFX1 U32(.A(flit42[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][32]));
	BUFX1 U33(.A(flit42[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][33]));
    NOR2X1 U34 ( .IN1(flit42[33]), .IN2(flit42[32]), .QN(norres_vc_buffer42_vc_buffer2) );
    OR4X1 U35 ( .IN1(flit42[29]), .IN2(flit42[28]), .IN3(flit42[27]), .IN4(flit42[26]), .Y(or1res_vc_buffer42) );
    OR4X1 U35 ( .IN1(flit42[25]), .IN2(flit42[24]), .IN3(flit42[23]), .IN4(flit42[22]), .Y(or2res_vc_buffer42) );
    OR2X1 U36 ( .A(or1res_vc_buffer42), .B(or2res_vc_buffer42), .Y(orres_vc_buffer42) );
    AND3X1 U37 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(norres_vc_buffer42_vc_buffer2), .IN3(orres_vc_buffer42), .Q(finres1_vc_buffer42) );
    MUX21X1 U38 (.IN1(next_locked_vc_buffer42), .IN2(1'b1), .S(finres1_vc_buffer42), .Q(next_locked_vc_buffer42);
    AND3X1 U39 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(flit42[33]), .IN3(flit42[32]), .Q(andres1_vc_buffer42) );
    MUX21X1 U40 (.IN1(next_locked_vc_buffer42), .IN2(1'b0), .S(andres1_vc_buffer42), .Q(next_locked_vc_buffer42);

    INVX1 U41 ( .A(full_vc_buffer42), .Y(full_vc_buffer42_not2) );
    INVX1 U42 ( .A(locked_by_route_ff_vc_buffer42), .Y(locked_by_route_ff_vc_buffer42_not2) );

    MUX21X1 U43 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer42_not2), .S(norres_vc_buffer42_vc_buffer2), .Q(thirdand_vc_buffer42);
    AND3X1 U44 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(full_vc_buffer42_not2), .IN3(thirdand_vc_buffer42), .Q(write_flit42_vc_buffer24) );
    AND2X1 U45 ( .IN1(full_vc_buffer42_not2), .IN2(norres_vc_buffer42_vc_buffer2), .Q(from_input_resp_input_datapath4[2]) );
    INVX1 U46 ( .A(empty_vc_buffer42), .Y(to_output_req_in_jump_input_datapath4put_datapath4[74]) );
    AND2X1 U47 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[74]), .IN2(to_output_resp_input_datapath4[2]), .Q(read_flit42_vc_buffer24) );
	BUFX1 U48(.A(to_output_req_in_jump_input_datapath4put_datapath4[76:75]), .Y(2'b10));

	DFFX2 U49 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U50 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U51 (.IN1(next_locked_vc_buffer42), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer42);

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath4put_datapath4[77]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath4put_datapath4[78]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath4put_datapath4[79]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath4put_datapath4[80]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath4put_datapath4[81]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath4put_datapath4[82]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath4put_datapath4[83]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath4put_datapath4[84]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath4put_datapath4[85]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath4put_datapath4[86]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath4put_datapath4[87]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath4put_datapath4[88]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath4put_datapath4[89]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath4put_datapath4[90]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath4put_datapath4[91]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath4put_datapath4[92]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath4put_datapath4[93]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath4put_datapath4[94]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath4put_datapath4[95]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath4put_datapath4[96]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath4put_datapath4[97]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath4put_datapath4[98]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath4put_datapath4[99]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath4put_datapath4[100]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath4put_datapath4[101]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath4put_datapath4[102]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath4put_datapath4[103]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath4put_datapath4[104]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath4put_datapath4[105]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath4put_datapath4[106]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath4put_datapath4[107]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath4put_datapath4[108]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath4put_datapath4[109]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath4put_datapath4[110]), .Y(ext_req_v_i[184:148][36]));
    XNOR2X1 U222 ( .IN1(ext_req_v_i[184:148][1]), .IN2(i_input_datapath4[0]), .QN(xnor1resu_input_datapath4) );
    XNOR2X1 U222 ( .IN1(ext_req_v_i[184:148][2]), .IN2(i_input_datapath4[1]), .QN(xnor2resu_input_datapath4) );
    AND2X1 U128 ( .IN1(xnor1resu_input_datapath4), .IN2(xnor2resu_input_datapath4), .Q(and1resu_input_datapath4) );
    AND3X1 U128 ( .IN1(and1resu_input_datapath4), .IN2(ext_req_v_i[184:148][0]), .IN2(ext_req_v_i[184:148][0]), .Q(cond1line_input_datapath4) );
    MUX21X1 U0009 (.IN1(vc_ch_act_in_input_datapath4[0]), .IN2(i_input_datapath4[0]), .S(cond1line_input_datapath4), .Q(vc_ch_act_in_input_datapath4[0]));
    MUX21X1 U0010 (.IN1(vc_ch_act_in_input_datapath4[1]), .IN2(i_input_datapath4[1]), .S(cond1line_input_datapath4), .Q(vc_ch_act_in_input_datapath4[1]));
    MUX21X1 U0011 (.IN1(req_in_jump_input_datapath4), .IN2(1), .S(cond1line_input_datapath4), .Q(req_in_jump_input_datapath4));
	BUFX1 U3(.A(from_input_req_in_jump_input_datapath4put_datapath4[40]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath4put_datapath4[41]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath4put_datapath4[42]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath4put_datapath4[43]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath4put_datapath4[44]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath4put_datapath4[45]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath4put_datapath4[46]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath4put_datapath4[47]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath4put_datapath4[48]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath4put_datapath4[49]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath4put_datapath4[50]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath4put_datapath4[51]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath4put_datapath4[52]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath4put_datapath4[53]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath4put_datapath4[54]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath4put_datapath4[55]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath4put_datapath4[56]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath4put_datapath4[57]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath4put_datapath4[58]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath4put_datapath4[59]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath4put_datapath4[60]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath4put_datapath4[61]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath4put_datapath4[62]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath4put_datapath4[63]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath4put_datapath4[64]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath4put_datapath4[65]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath4put_datapath4[66]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath4put_datapath4[67]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath4put_datapath4[68]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath4put_datapath4[69]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath4put_datapath4[70]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath4put_datapath4[71]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath4put_datapath4[72]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath4put_datapath4[73]), .Y(ext_req_v_i[184:148][36]));

	BUFX1 U3(.A(from_input_req_in_jump_input_datapath4put_datapath4[3]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U4(.A(from_input_req_in_jump_input_datapath4put_datapath4[4]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U5(.A(from_input_req_in_jump_input_datapath4put_datapath4[5]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U6(.A(from_input_req_in_jump_input_datapath4put_datapath4[6]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U7(.A(from_input_req_in_jump_input_datapath4put_datapath4[7]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U8(.A(from_input_req_in_jump_input_datapath4put_datapath4[8]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U9(.A(from_input_req_in_jump_input_datapath4put_datapath4[9]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U10(.A(from_input_req_in_jump_input_datapath4put_datapath4[10]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U11(.A(from_input_req_in_jump_input_datapath4put_datapath4[11]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U12(.A(from_input_req_in_jump_input_datapath4put_datapath4[12]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U13(.A(from_input_req_in_jump_input_datapath4put_datapath4[13]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U14(.A(from_input_req_in_jump_input_datapath4put_datapath4[14]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U15(.A(from_input_req_in_jump_input_datapath4put_datapath4[15]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U16(.A(from_input_req_in_jump_input_datapath4put_datapath4[16]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U17(.A(from_input_req_in_jump_input_datapath4put_datapath4[17]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U18(.A(from_input_req_in_jump_input_datapath4put_datapath4[18]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U19(.A(from_input_req_in_jump_input_datapath4put_datapath4[19]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U20(.A(from_input_req_in_jump_input_datapath4put_datapath4[20]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U21(.A(from_input_req_in_jump_input_datapath4put_datapath4[21]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U22(.A(from_input_req_in_jump_input_datapath4put_datapath4[22]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U23(.A(from_input_req_in_jump_input_datapath4put_datapath4[23]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U24(.A(from_input_req_in_jump_input_datapath4put_datapath4[24]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U25(.A(from_input_req_in_jump_input_datapath4put_datapath4[25]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U26(.A(from_input_req_in_jump_input_datapath4put_datapath4[26]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U27(.A(from_input_req_in_jump_input_datapath4put_datapath4[27]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U28(.A(from_input_req_in_jump_input_datapath4put_datapath4[28]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U29(.A(from_input_req_in_jump_input_datapath4put_datapath4[29]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U30(.A(from_input_req_in_jump_input_datapath4put_datapath4[30]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U31(.A(from_input_req_in_jump_input_datapath4put_datapath4[31]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U32(.A(from_input_req_in_jump_input_datapath4put_datapath4[32]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U33(.A(from_input_req_in_jump_input_datapath4put_datapath4[33]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U34(.A(from_input_req_in_jump_input_datapath4put_datapath4[34]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U35(.A(from_input_req_in_jump_input_datapath4put_datapath4[35]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U36(.A(from_input_req_in_jump_input_datapath4put_datapath4[36]), .Y(ext_req_v_i[184:148][36]));

    MUX21X1 U0012 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4 * 37]), .IN2(ext_req_v_i[184:148][0]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4 * 37]));
    MUX21X1 U0013 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+2]), .IN2(vc_ch_act_in_input_datapath4[1]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+2]));
    MUX21X1 U0014 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+1]), .IN2(vc_ch_act_in_input_datapath4[0]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+1]));
    MUX21X1 U0015 (.IN1(ext_resp_v_o[5:4][0]), .IN2(from_input_resp_input_datapath4[vc_ch_act_in_input_datapath4]), .S(req_in_jump_input_datapath4), .Q(ext_resp_v_o[5:4][0]));

    INVX1 U041 ( .A(req_in_jump_input_datapath4), .Y(req_in_jump_input_datapath4_not) );
    MUX21X1 U0016 (.IN1(ext_resp_v_o[5:4][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath4_not), .Q(ext_resp_v_o[5:4][0]));
    BUFX1 U34(.A(from_input_req_in_jump_input_datapath4put_datapath4[34]), .Y(ext_req_v_i[184:148][34]));

    XOR2X1 U0222 ( .IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b1), .Q(xor1resu_input_datapath4) );
    MUX21X1 U0017 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(xor1resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U0018 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b0), .S(xor1resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[1]));
    AND2X1 U38123 ( .IN1(xor1resu_input_datapath4), .IN2(to_output_req_in_jump_input_datapath4put_datapath4[j_input_datapath4*37]), .Q(and2resu_input_datapath4) );
    MUX21X1 U0019 (.IN1(vc_ch_act_out_input_datapath4[0]), .IN2(j_input_datapath4[0]), .S(and2resu_input_datapath4), .Q(vc_ch_act_out_input_datapath4[0]));
    MUX21X1 U0020 (.IN1(vc_ch_act_out_input_datapath4[1]), .IN2(j_input_datapath4[1]), .S(and2resu_input_datapath4), .Q(vc_ch_act_out_input_datapath4[1]));
    MUX21X1 U0021 (.IN1(req_out_jump_input_datapath4), .IN2(1'b1), .S(and2resu_input_datapath4), .Q(req_out_jump_input_datapath4));
    MUX21X1 U0022 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(and2resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U0023 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b1), .S(and2resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[1]));
    HADDX1 U00021 ( .A0(j_input_datapath4[0]), .B0(1'b1), .C1(j_input_datapath4[1]), .SO(j_input_datapath4[0]) );
    HADDX1 U00022 ( .A0(j_input_datapath4[0]), .B0(1'b1), .C1(j_input_datapath4[1]), .SO(j_input_datapath4[0]) );
    AND2X1 U38111 ( .IN1(xor1resu_input_datapath4), .IN2(to_output_req_in_jump_input_datapath4put_datapath4[j_input_datapath4*37]), .Q(and3resu) );
    NAND2X1 U29311(.A(_sv2v_jump_input_datapath4[0]),.B(_sv2v_jump_input_datapath4[1]),.Y(nand1resu_input_datapath44));
    MUX21X1 U00212 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(nand1resu_input_datapath44), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U00213 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b0), .S(nand1resu_input_datapath44), .Q(_sv2v_jump_input_datapath4[1]));
    XNOR2X1 U17581 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(_sv2v_jump_input_datapath4[1]), .Q(xnor23resu_input_datapath4) );
    AND2X1 U38111 ( .IN1(xnor23resu_input_datapath4), .IN2(req_out_jump_input_datapath4), .Q(and4resu_input_datapath4) );

    MUX21X1 U3(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[184:148][3]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U4(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[184:148][4]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U5(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[184:148][5]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U6(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[184:148][6]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U7(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[184:148][7]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U8(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[184:148][8]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U9(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[184:148][9]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U10(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[184:148][10]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U11(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[184:148][11]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U12(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[184:148][12]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U13(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[184:148][13]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U14(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[184:148][14]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U15(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[184:148][15]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U16(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[184:148][16]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U17(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[184:148][17]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U18(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[184:148][18]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U19(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[184:148][19]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U20(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[184:148][20]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U21(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[184:148][21]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U22(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[184:148][22]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U23(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[184:148][23]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U24(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[184:148][24]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U25(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[184:148][25]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U26(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[184:148][26]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U27(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[184:148][27]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U28(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[184:148][28]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U29(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[184:148][29]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U30(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[184:148][30]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U31(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[184:148][31]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U32(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[184:148][32]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U33(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[184:148][33]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U34(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[184:148][34]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U35(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[184:148][35]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U36(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[184:148][36]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U321111(.IN1(int_req_v[184:148][0]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4 * 37)]), .S(and4resu_input_datapath4), .Q(int_req_v[184:148][0]));
	MUX21X1 U331112(.IN1(int_req_v[184:148][1]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+1]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+1]));
	MUX21X1 U331122(.IN1(int_req_v[184:148][2]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+2]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+2]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4]),.IN2(int_resp_v[5:4]), .S(and4resu_input_datapath4), .Q(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4]));
	MUX21X1 U352221(.IN1(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4+1]),.IN2(int_resp_v[5:4]), .S(and4resu_input_datapath4), .Q(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4+1]));



//output part	

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1[0]), .Y(i_0_not_high_prior_arbiter1) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1[0]), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(_sv2v_jump_high_prior_arbiter1[1]), .QN(nandres_high_prior_arbiter1) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2[0]), .Y(i_0_not_high_prior_arbiter2) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2[0]), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(_sv2v_jump_high_prior_arbiter2[1]), .QN(nandres_high_prior_arbiter2) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter[0]), .B(valid_from_im_output_module[3:0][0]), .Y(mask_req_rr_arbiter[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter[1]), .B(valid_from_im_output_module[3:0][1]), .Y(mask_req_rr_arbiter[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter[0]), .Y(next_mask_rr_arbiter[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter[1]), .Y(next_mask_rr_arbiter[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter[0]), .IN2(raw_grant_rr_arbiter[0]), .S(xnor0res_rr_arbiter), .Q(grant_im_output_module[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter[1]), .IN2(raw_grant_rr_arbiter[1]), .S(xnor1res_rr_arbiter), .Q(grant_im_output_module[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter[1]), .B(1'b0), .Y(firstif_rr_arbiter) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter), .B(grant_im_output_module[3:0][i_rr_arbiter[0]]), .Y(secondif_rr_arbiter) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[1]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter[0]), .Q(j_rr_arbiter[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter), .B(j_rr_arbiter[0]), .Y(thirdif_rr_arbiter) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter[j_rr_arbiter[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter), .Q(next_mask_rr_arbiter[j_rr_arbiter[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b1), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(_sv2v_jump_rr_rr_arbiter[1]), .QN(fourthif_rr_arbiter) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter[0]), .IN2(next_mask_rr_arbiter[0]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter[1]), .IN2(next_mask_rr_arbiter[1]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter), .IN2(1'sb1), .S(arst_value_rr_arbiter), .Q(mask_ff_rr_arbiter[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter11) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter11[0]), .Y(i_0_not_high_prior_arbiter11) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter11), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter11[0]), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b1), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(_sv2v_jump_high_prior_arbiter11[1]), .QN(nandres_high_prior_arbiter11) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter21[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter21[0]), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(_sv2v_jump_high_prior_arbiter21[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter1[0]), .B(valid_from_im_output_module[7:4][0]), .Y(mask_req_rr_arbiter1[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter1[1]), .B(valid_from_im_output_module[7:4][1]), .Y(mask_req_rr_arbiter1[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter1[0]), .Y(next_mask_rr_arbiter1[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter1[1]), .Y(next_mask_rr_arbiter1[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter1[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter1) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter1[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter1) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter1[0]), .IN2(raw_grant_rr_arbiter1[0]), .S(xnor0res_rr_arbiter1), .Q(grant_im_output_module[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter1[1]), .IN2(raw_grant_rr_arbiter1[1]), .S(xnor1res_rr_arbiter1), .Q(grant_im_output_module[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter1[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter1[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter1[1]), .B(1'b0), .Y(firstif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter1), .B(grant_im_output_module[7:4][i_rr_arbiter1[0]]), .Y(secondif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[1]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter1[0]), .Q(j_rr_arbiter1[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter1), .B(j_rr_arbiter1[0]), .Y(thirdif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter1[j_rr_arbiter1[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter1), .Q(next_mask_rr_arbiter1[j_rr_arbiter1[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b1), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(_sv2v_jump_rr_rr_arbiter1[1]), .QN(fourthif_rr_arbiter1) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter1) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter1) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter1[0]), .IN2(next_mask_rr_arbiter1[0]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter1[1]), .IN2(next_mask_rr_arbiter1[1]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter11), .IN2(1'sb1), .S(arst_value_rr_arbiter1), .Q(mask_ff_rr_arbiter1[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter12) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter12[0]), .Y(i_0_not_high_prior_arbiter12) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter12), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter12[0]), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b1), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(_sv2v_jump_high_prior_arbiter12[1]), .QN(nandres_high_prior_arbiter12) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter22[0]), .Y(i_0_not_high_prior_arbiter22) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter22[0]), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(_sv2v_jump_high_prior_arbiter22[1]), .QN(nandres_high_prior_arbiter22) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter2[0]), .B(valid_from_im_output_module[11:8][0]), .Y(mask_req_rr_arbiter2[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter2[1]), .B(valid_from_im_output_module[11:8][1]), .Y(mask_req_rr_arbiter2[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter2[0]), .Y(next_mask_rr_arbiter2[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter2[1]), .Y(next_mask_rr_arbiter2[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter2[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter2) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter2[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter2) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter2[0]), .IN2(raw_grant_rr_arbiter2[0]), .S(xnor0res_rr_arbiter2), .Q(grant_im_output_module[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter2[1]), .IN2(raw_grant_rr_arbiter2[1]), .S(xnor1res_rr_arbiter2), .Q(grant_im_output_module[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter2[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter2[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter2[1]), .B(1'b0), .Y(firstif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter2), .B(grant_im_output_module[11:8][i_rr_arbiter2[0]]), .Y(secondif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[1]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter2[0]), .Q(j_rr_arbiter2[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter2), .B(j_rr_arbiter2[0]), .Y(thirdif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter2[j_rr_arbiter2[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter2), .Q(next_mask_rr_arbiter2[j_rr_arbiter2[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b1), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(_sv2v_jump_rr_rr_arbiter2[1]), .QN(fourthif_rr_arbiter2) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter2) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter2) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter2[0]), .IN2(next_mask_rr_arbiter2[0]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter2[1]), .IN2(next_mask_rr_arbiter2[1]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter22), .IN2(1'sb1), .S(arst_value_rr_arbiter2), .Q(mask_ff_rr_arbiter2[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37]), .IN2(vc_channel_output_module[1]), .QN(xnor1resu1_output_module) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37-1]), .IN2(vc_channel_output_module[0]), .QN(xnor2resu1_output_module) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module), .IN2(xnor2resu1_output_module), .Q(and1resu1_output_module) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]), .IN2(1'b1), .S(and1resu1_output_module), .Q(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .Q(xor1resu1_output_module) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module_1[0]), .IN2(_sv2v_jump_output_module[0]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module_1[1]), .IN2(_sv2v_jump_output_module[1]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[vc_channel_output_module[1:0]*4+in_mod_output_module[1:0]]), .Q(and2resu1_output_module) );

    MUX21X1 U3(.IN1(head_flit_output_module[3]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+3]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[3]));
	MUX21X1 U4(.IN1(head_flit_output_module[4]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+4]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[4]));
	MUX21X1 U5(.IN1(head_flit_output_module[5]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+5]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[5]));
	MUX21X1 U6(.IN1(head_flit_output_module[6]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+6]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[6]));
	MUX21X1 U7(.IN1(head_flit_output_module[7]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+7]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[7]));
	MUX21X1 U8(.IN1(head_flit_output_module[8]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+8]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[8]));
	MUX21X1 U9(.IN1(head_flit_output_module[9]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+9]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[9]));
	MUX21X1 U10(.IN1(head_flit_output_module[10]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+10]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[10]));
	MUX21X1 U11(.IN1(head_flit_output_module[11]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+11]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[11]));
	MUX21X1 U12(.IN1(head_flit_output_module[12]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+12]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[12]));
	MUX21X1 U13(.IN1(head_flit_output_module[13]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+13]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[13]));
	MUX21X1 U14(.IN1(head_flit_output_module[14]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+14]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[14]));
	MUX21X1 U15(.IN1(head_flit_output_module[15]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+15]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[15]));
	MUX21X1 U16(.IN1(head_flit_output_module[16]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+16]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[16]));
	MUX21X1 U17(.IN1(head_flit_output_module[17]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+17]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[17]));
	MUX21X1 U18(.IN1(head_flit_output_module[18]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+18]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[18]));
	MUX21X1 U19(.IN1(head_flit_output_module[19]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+19]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[19]));
	MUX21X1 U20(.IN1(head_flit_output_module[20]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+20]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[20]));
	MUX21X1 U21(.IN1(head_flit_output_module[21]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+21]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[21]));
	MUX21X1 U22(.IN1(head_flit_output_module[22]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+22]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[22]));
	MUX21X1 U23(.IN1(head_flit_output_module[23]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+23]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[23]));
	MUX21X1 U24(.IN1(head_flit_output_module[24]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+24]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[24]));
	MUX21X1 U25(.IN1(head_flit_output_module[25]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+25]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[25]));
	MUX21X1 U26(.IN1(head_flit_output_module[26]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+26]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[26]));
	MUX21X1 U27(.IN1(head_flit_output_module[27]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+27]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[27]));
	MUX21X1 U28(.IN1(head_flit_output_module[28]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+28]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[28]));
	MUX21X1 U29(.IN1(head_flit_output_module[29]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+29]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[29]));
	MUX21X1 U30(.IN1(head_flit_output_module[30]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+30]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[30]));
	MUX21X1 U31(.IN1(head_flit_output_module[31]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+31]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[31]));
	MUX21X1 U32(.IN1(head_flit_output_module[32]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+32]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[32]));
	MUX21X1 U33(.IN1(head_flit_output_module[33]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+33]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[33]));
	MUX21X1 U34(.IN1(head_flit_output_module[34]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+34]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[34]));
	MUX21X1 U35(.IN1(head_flit_output_module[35]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+35]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[35]));
	MUX21X1 U36(.IN1(head_flit_output_module[36]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+36]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[36]));

    INVX1 U041 ( .A(head_flit_output_module[32]), .Y(head_flit_output_module_32_not_output_module) );
    AND2X1 U1218 ( .IN1(head_flit_output_module_32_not_output_module), .IN2(head_flit_output_module[33]), .Q(and3resu1_output_module) );
    NOR4X1 U175821 (.IN1(head_flit_output_module[29]), .IN2(head_flit_output_module[28]), .IN3(head_flit_output_module[27]), .IN4(head_flit_output_module[26]), .Q(nor23resu1_output_module) );
    NOR4X1 U175831 (.IN1(head_flit_output_module[25]), .IN2(head_flit_output_module[24]), .IN3(head_flit_output_module[23]), .IN4(head_flit_output_module[22]), .Q(nor23resu2_output_module) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module), .IN2(nor23resu2_output_module), .Q(and4resu1_output_module) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module[33]), .IN2(head_flit_output_module[32]), .Q(nor23resu3_output_module) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module), .IN2(and4resu1_output_module), .Q(and5resu1_output_module) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module), .IN2(nor23resu3_output_module), .Q(or12resu12_output_module) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[1:0][0]), .IN2(or12resu12_output_module), .Q(and6resu1_output_module) );    
	MUX21X1 U361(.IN1(tail_flit_im_output_module[vc_channel_output_module[1:0]]), .IN2(and6resu1_output_module), .S(and2resu1_output_module) ,.Q(tail_flit_im_output_module[vc_channel_output_module[1:0]]);
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module[0]),.B(_sv2v_jump_output_module[1]),.Y(nand1resu_output_module));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module), .IN2(nand1resu_output_module), .Q(and7resu1) );    
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(_sv2v_jump_output_module_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U00021 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );



	BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module[0]));
	BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[i_output_module[1:0] * 4+:4]), .Q(and8resu1_output_module) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module[0]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[0]);
	MUX21X1 U3631(.IN1(vc_ch_act_out_output_module[1]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[1]);
	MUX21X1 U3631(.IN1(req_out_output_module), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(req_out_output_module);
	MUX21X1 U3621(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3631(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module[1]), .Q(norfinresu1_output_module) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module), .IN2(req_out_output_module), .Q(and9resu1_output_module) );    
	HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module), .IN2(grant_im_output_module[(vc_ch_act_out_output_module * 4) + i_output_module[1:0]]), .Q(and10resu1_output_module) );    

	MUX21X1 U3(.IN1(ext_req_v_o[36:0][3]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+3]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][3]));
	MUX21X1 U4(.IN1(ext_req_v_o[36:0][4]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+4]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][4]));
	MUX21X1 U5(.IN1(ext_req_v_o[36:0][5]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+5]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][5]));
	MUX21X1 U6(.IN1(ext_req_v_o[36:0][6]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+6]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][6]));
	MUX21X1 U7(.IN1(ext_req_v_o[36:0][7]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+7]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][7]));
	MUX21X1 U8(.IN1(ext_req_v_o[36:0][8]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+8]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][8]));
	MUX21X1 U9(.IN1(ext_req_v_o[36:0][9]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+9]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][9]));
	MUX21X1 U10(.IN1(ext_req_v_o[36:0][10]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+10]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][10]));
	MUX21X1 U11(.IN1(ext_req_v_o[36:0][11]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+11]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][11]));
	MUX21X1 U12(.IN1(ext_req_v_o[36:0][12]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+12]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][12]));
	MUX21X1 U13(.IN1(ext_req_v_o[36:0][13]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+13]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][13]));
	MUX21X1 U14(.IN1(ext_req_v_o[36:0][14]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+14]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][14]));
	MUX21X1 U15(.IN1(ext_req_v_o[36:0][15]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+15]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][15]));
	MUX21X1 U16(.IN1(ext_req_v_o[36:0][16]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+16]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][16]));
	MUX21X1 U17(.IN1(ext_req_v_o[36:0][17]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+17]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][17]));
	MUX21X1 U18(.IN1(ext_req_v_o[36:0][18]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+18]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][18]));
	MUX21X1 U19(.IN1(ext_req_v_o[36:0][19]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+19]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][19]));
	MUX21X1 U20(.IN1(ext_req_v_o[36:0][20]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+20]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][20]));
	MUX21X1 U21(.IN1(ext_req_v_o[36:0][21]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+21]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][21]));
	MUX21X1 U22(.IN1(ext_req_v_o[36:0][22]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+22]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][22]));
	MUX21X1 U23(.IN1(ext_req_v_o[36:0][23]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+23]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][23]));
	MUX21X1 U24(.IN1(ext_req_v_o[36:0][24]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+24]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][24]));
	MUX21X1 U25(.IN1(ext_req_v_o[36:0][25]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+25]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][25]));
	MUX21X1 U26(.IN1(ext_req_v_o[36:0][26]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+26]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][26]));
	MUX21X1 U27(.IN1(ext_req_v_o[36:0][27]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+27]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][27]));
	MUX21X1 U28(.IN1(ext_req_v_o[36:0][28]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+28]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][28]));
	MUX21X1 U29(.IN1(ext_req_v_o[36:0][29]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+29]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][29]));
	MUX21X1 U30(.IN1(ext_req_v_o[36:0][30]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+30]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][30]));
	MUX21X1 U31(.IN1(ext_req_v_o[36:0][31]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+31]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][31]));
	MUX21X1 U32(.IN1(ext_req_v_o[36:0][32]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+32]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][32]));
	MUX21X1 U33(.IN1(ext_req_v_o[36:0][33]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+33]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][33]));
	MUX21X1 U34(.IN1(ext_req_v_o[36:0][34]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+34]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][34]));
	MUX21X1 U35(.IN1(ext_req_v_o[36:0][35]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+35]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][35]));
	MUX21X1 U36(.IN1(ext_req_v_o[36:0][36]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+36]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][36]));

	MUX21X1 U36221(.IN1(ext_req_v_o[36:0][0]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][0]);
	MUX21X1 U36221(.IN1(ext_req_v_o[36:0][1]), .IN2(vc_ch_act_out_output_module[0]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][1]);
	MUX21X1 U36331(.IN1(ext_req_v_o[36:0][2]), .IN2(vc_ch_act_out_output_module[1]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][2]);    
	MUX21X1 U36221(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U36331(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module), .IN2(nand1resu_output_module), .Q(and11resu1_output_module) );    
	MUX21X1 U36221(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U36331(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);  





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter111[0]), .Y(i_0_not_high_prior_arbiter111) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter111), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter111[0]), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(_sv2v_jump_high_prior_arbiter111[1]), .QN(nandres_high_prior_arbiter111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter211[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter211[0]), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(_sv2v_jump_high_prior_arbiter211[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter11[0]), .B(valid_from_im_output_module1[3:0][0]), .Y(mask_req_rr_arbiter11[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter11[1]), .B(valid_from_im_output_module1[3:0][1]), .Y(mask_req_rr_arbiter11[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter11[0]), .Y(next_mask_rr_arbiter11[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter11[1]), .Y(next_mask_rr_arbiter11[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter11[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter11) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter11[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter11) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter11[0]), .IN2(raw_grant_rr_arbiter11[0]), .S(xnor0res_rr_arbiter11), .Q(grant_im_output_module1[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter11[1]), .IN2(raw_grant_rr_arbiter11[1]), .S(xnor1res_rr_arbiter11), .Q(grant_im_output_module1[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter11[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter11[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter11[1]), .B(1'b0), .Y(firstif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter11), .B(grant_im_output_module1[3:0][i_rr_arbiter11[0]]), .Y(secondif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[1]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter11[0]), .Q(j_rr_arbiter11[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter11), .B(j_rr_arbiter11[0]), .Y(thirdif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter11[j_rr_arbiter11[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter11), .Q(next_mask_rr_arbiter11[j_rr_arbiter11[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b1), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(_sv2v_jump_rr_rr_arbiter11[1]), .QN(fourthif_rr_arbiter11) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter11) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter11) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter11[0]), .IN2(next_mask_rr_arbiter11[0]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter11[1]), .IN2(next_mask_rr_arbiter11[1]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter1111), .IN2(1'sb1), .S(arst_value_rr_arbiter11), .Q(mask_ff_rr_arbiter11[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1111[0]), .Y(i_0_not_high_prior_arbiter1111) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1111), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1111[0]), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(_sv2v_jump_high_prior_arbiter1111[1]), .QN(nandres_high_prior_arbiter1111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2111) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2111[0]), .Y(i_0_not_high_prior_arbiter2111) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2111), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2111[0]), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(_sv2v_jump_high_prior_arbiter2111[1]), .QN(nandres_high_prior_arbiter2111) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter111[0]), .B(valid_from_im_output_module1[7:4][0]), .Y(mask_req_rr_arbiter111[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter111[1]), .B(valid_from_im_output_module1[7:4][1]), .Y(mask_req_rr_arbiter111[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter111[0]), .Y(next_mask_rr_arbiter111[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter111[1]), .Y(next_mask_rr_arbiter111[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter111[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter111) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter111[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter111) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter111[0]), .IN2(raw_grant_rr_arbiter111[0]), .S(xnor0res_rr_arbiter111), .Q(grant_im_output_module1[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter111[1]), .IN2(raw_grant_rr_arbiter111[1]), .S(xnor1res_rr_arbiter111), .Q(grant_im_output_module1[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter111[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter111[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter111[1]), .B(1'b0), .Y(firstif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter111), .B(grant_im_output_module1[7:4][i_rr_arbiter111[0]]), .Y(secondif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[1]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter111[0]), .Q(j_rr_arbiter111[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter111), .B(j_rr_arbiter111[0]), .Y(thirdif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter111[j_rr_arbiter111[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter111), .Q(next_mask_rr_arbiter111[j_rr_arbiter111[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b1), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(_sv2v_jump_rr_rr_arbiter111[1]), .QN(fourthif_rr_arbiter111) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter111) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter111) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter111[0]), .IN2(next_mask_rr_arbiter111[0]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter111[1]), .IN2(next_mask_rr_arbiter111[1]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter111111), .IN2(1'sb1), .S(arst_value_rr_arbiter111), .Q(mask_ff_rr_arbiter111[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1112) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1112[0]), .Y(i_0_not_high_prior_arbiter1112) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1112), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1112[0]), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b1), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(_sv2v_jump_high_prior_arbiter1112[1]), .QN(nandres_high_prior_arbiter1112) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter212) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2112[0]), .Y(i_0_not_high_prior_arbiter212) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter212), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2112[0]), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(_sv2v_jump_high_prior_arbiter2112[1]), .QN(nandres_high_prior_arbiter212) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter112[0]), .B(valid_from_im_output_module1[11:8][0]), .Y(mask_req_rr_arbiter112[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter112[1]), .B(valid_from_im_output_module1[11:8][1]), .Y(mask_req_rr_arbiter112[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter112[0]), .Y(next_mask_rr_arbiter112[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter112[1]), .Y(next_mask_rr_arbiter112[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter112[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter112) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter112[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter112) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter112[0]), .IN2(raw_grant_rr_arbiter112[0]), .S(xnor0res_rr_arbiter112), .Q(grant_im_output_module1[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter112[1]), .IN2(raw_grant_rr_arbiter112[1]), .S(xnor1res_rr_arbiter112), .Q(grant_im_output_module1[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter112[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter112[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter112[1]), .B(1'b0), .Y(firstif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter112), .B(grant_im_output_module1[11:8][i_rr_arbiter112[0]]), .Y(secondif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[1]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter112[0]), .Q(j_rr_arbiter112[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter112), .B(j_rr_arbiter112[0]), .Y(thirdif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter112[j_rr_arbiter112[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter112), .Q(next_mask_rr_arbiter112[j_rr_arbiter112[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b1), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(_sv2v_jump_rr_rr_arbiter112[1]), .QN(fourthif_rr_arbiter112) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter112) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter112) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter112[0]), .IN2(next_mask_rr_arbiter112[0]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter112[1]), .IN2(next_mask_rr_arbiter112[1]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter111122), .IN2(1'sb1), .S(arst_value_rr_arbiter112), .Q(mask_ff_rr_arbiter112[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37]), .IN2(vc_channel_output_module1[1]), .QN(xnor1resu1_output_module1) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37-1]), .IN2(vc_channel_output_module1[0]), .QN(xnor2resu1_output_module1) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module1), .IN2(xnor2resu1_output_module1), .Q(and1resu1_output_module1) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]), .IN2(1'b1), .S(and1resu1_output_module1), .Q(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .Q(xor1resu1_output_module1) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module1_1[0]), .IN2(_sv2v_jump_output_module1[0]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module1_1[1]), .IN2(_sv2v_jump_output_module1[1]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[vc_channel_output_module1[1:0]*4+in_mod_output_module1[1:0]]), .Q(and2resu1_output_module1) );

    MUX21X1 U3(.IN1(head_flit_output_module1[3]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+3]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[3]));
    MUX21X1 U4(.IN1(head_flit_output_module1[4]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+4]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[4]));
    MUX21X1 U5(.IN1(head_flit_output_module1[5]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+5]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[5]));
    MUX21X1 U6(.IN1(head_flit_output_module1[6]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+6]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[6]));
    MUX21X1 U7(.IN1(head_flit_output_module1[7]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+7]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[7]));
    MUX21X1 U8(.IN1(head_flit_output_module1[8]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+8]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[8]));
    MUX21X1 U9(.IN1(head_flit_output_module1[9]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+9]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[9]));
    MUX21X1 U10(.IN1(head_flit_output_module1[10]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+10]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[10]));
    MUX21X1 U11(.IN1(head_flit_output_module1[11]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+11]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[11]));
    MUX21X1 U12(.IN1(head_flit_output_module1[12]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+12]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[12]));
    MUX21X1 U13(.IN1(head_flit_output_module1[13]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+13]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[13]));
    MUX21X1 U14(.IN1(head_flit_output_module1[14]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+14]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[14]));
    MUX21X1 U15(.IN1(head_flit_output_module1[15]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+15]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[15]));
    MUX21X1 U16(.IN1(head_flit_output_module1[16]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+16]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[16]));
    MUX21X1 U17(.IN1(head_flit_output_module1[17]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+17]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[17]));
    MUX21X1 U18(.IN1(head_flit_output_module1[18]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+18]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[18]));
    MUX21X1 U19(.IN1(head_flit_output_module1[19]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+19]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[19]));
    MUX21X1 U20(.IN1(head_flit_output_module1[20]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+20]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[20]));
    MUX21X1 U21(.IN1(head_flit_output_module1[21]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+21]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[21]));
    MUX21X1 U22(.IN1(head_flit_output_module1[22]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+22]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[22]));
    MUX21X1 U23(.IN1(head_flit_output_module1[23]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+23]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[23]));
    MUX21X1 U24(.IN1(head_flit_output_module1[24]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+24]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[24]));
    MUX21X1 U25(.IN1(head_flit_output_module1[25]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+25]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[25]));
    MUX21X1 U26(.IN1(head_flit_output_module1[26]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+26]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[26]));
    MUX21X1 U27(.IN1(head_flit_output_module1[27]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+27]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[27]));
    MUX21X1 U28(.IN1(head_flit_output_module1[28]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+28]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[28]));
    MUX21X1 U29(.IN1(head_flit_output_module1[29]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+29]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[29]));
    MUX21X1 U30(.IN1(head_flit_output_module1[30]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+30]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[30]));
    MUX21X1 U31(.IN1(head_flit_output_module1[31]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+31]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[31]));
    MUX21X1 U32(.IN1(head_flit_output_module1[32]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+32]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[32]));
    MUX21X1 U33(.IN1(head_flit_output_module1[33]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+33]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[33]));
    MUX21X1 U34(.IN1(head_flit_output_module1[34]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+34]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[34]));
    MUX21X1 U35(.IN1(head_flit_output_module1[35]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+35]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[35]));
    MUX21X1 U36(.IN1(head_flit_output_module1[36]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+36]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[36]));

    INVX1 U041 ( .A(head_flit_output_module1[32]), .Y(head_flit_output_module1_32_not_output_module1) );
    AND2X1 U1218 ( .IN1(head_flit_output_module1_32_not_output_module1), .IN2(head_flit_output_module1[33]), .Q(and3resu1_output_module1) );
    NOR4X1 U175821 (.IN1(head_flit_output_module1[29]), .IN2(head_flit_output_module1[28]), .IN3(head_flit_output_module1[27]), .IN4(head_flit_output_module1[26]), .Q(nor23resu1_output_module1) );
    NOR4X1 U175831 (.IN1(head_flit_output_module1[25]), .IN2(head_flit_output_module1[24]), .IN3(head_flit_output_module1[23]), .IN4(head_flit_output_module1[22]), .Q(nor23resu2_output_module1) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module1), .IN2(nor23resu2_output_module1), .Q(and4resu1_output_module1) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module1[33]), .IN2(head_flit_output_module1[32]), .Q(nor23resu3_output_module1) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module1), .IN2(and4resu1_output_module1), .Q(and5resu1_output_module1) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module1), .IN2(nor23resu3_output_module1), .Q(or12resu12_output_module1) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[2:1][0]), .IN2(or12resu12_output_module1), .Q(and6resu1_output_module1) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]), .IN2(and6resu1_output_module1), .S(and2resu1_output_module1) ,.Q(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module1[0]),.B(_sv2v_jump_output_module1[1]),.Y(nand1resu_output_module1));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(_sv2v_jump_output_module1_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module1[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module1[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[i_output_module1[1:0] * 4+:4]), .Q(and8resu1_output_module1) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module1[0]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module1[1]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[1]);
    MUX21X1 U3631(.IN1(req_out_output_module1), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(req_out_output_module1);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1[1]), .Q(norfinresu1_output_module1) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module1), .IN2(req_out_output_module1), .Q(and9resu1_output_module1) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module1), .IN2(grant_im_output_module1[(vc_ch_act_out_output_module1 * 4) + i_output_module1[1:0]]), .Q(and10resu1_output_module1) );    

    MUX21X1 U3(.IN1(ext_req_v_o[73:37][3]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+3]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[73:37][4]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+4]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[73:37][5]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+5]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[73:37][6]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+6]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[73:37][7]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+7]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[73:37][8]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+8]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[73:37][9]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+9]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[73:37][10]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+10]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[73:37][11]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+11]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[73:37][12]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+12]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[73:37][13]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+13]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[73:37][14]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+14]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[73:37][15]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+15]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[73:37][16]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+16]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[73:37][17]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+17]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[73:37][18]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+18]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[73:37][19]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+19]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[73:37][20]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+20]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[73:37][21]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+21]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[73:37][22]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+22]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[73:37][23]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+23]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[73:37][24]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+24]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[73:37][25]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+25]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[73:37][26]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+26]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[73:37][27]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+27]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[73:37][28]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+28]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[73:37][29]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+29]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[73:37][30]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+30]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[73:37][31]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+31]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[73:37][32]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+32]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[73:37][33]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+33]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[73:37][34]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+34]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[73:37][35]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+35]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[73:37][36]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+36]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[73:37][0]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[73:37][1]), .IN2(vc_ch_act_out_output_module1[0]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[73:37][2]), .IN2(vc_ch_act_out_output_module1[1]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and11resu1_output_module1) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    
    
 





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter122) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter122[0]), .Y(i_0_not_high_prior_arbiter122) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter122), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter122[0]), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b1), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(_sv2v_jump_high_prior_arbiter122[1]), .QN(nandres_high_prior_arbiter122) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter222[0]), .Y(i_0_not_high_prior_arbiter222) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter222), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter222[0]), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(_sv2v_jump_high_prior_arbiter222[1]), .QN(nandres_high_prior_arbiter222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter22[0]), .B(valid_from_im_output_module2[3:0][0]), .Y(mask_req_rr_arbiter22[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter22[1]), .B(valid_from_im_output_module2[3:0][1]), .Y(mask_req_rr_arbiter22[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter22[0]), .Y(next_mask_rr_arbiter22[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter22[1]), .Y(next_mask_rr_arbiter22[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter22[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter22) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter22[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter22) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter22[0]), .IN2(raw_grant_rr_arbiter22[0]), .S(xnor0res_rr_arbiter22), .Q(grant_im_output_module2[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter22[1]), .IN2(raw_grant_rr_arbiter22[1]), .S(xnor1res_rr_arbiter22), .Q(grant_im_output_module2[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter22[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter22[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter22[1]), .B(1'b0), .Y(firstif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter22), .B(grant_im_output_module2[3:0][i_rr_arbiter22[0]]), .Y(secondif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[1]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter22[0]), .Q(j_rr_arbiter22[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter22), .B(j_rr_arbiter22[0]), .Y(thirdif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter22[j_rr_arbiter22[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter22), .Q(next_mask_rr_arbiter22[j_rr_arbiter22[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b1), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(_sv2v_jump_rr_rr_arbiter22[1]), .QN(fourthif_rr_arbiter22) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter22) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter22) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter22[0]), .IN2(next_mask_rr_arbiter22[0]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter22[1]), .IN2(next_mask_rr_arbiter22[1]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter2222), .IN2(1'sb1), .S(arst_value_rr_arbiter22), .Q(mask_ff_rr_arbiter22[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1221) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1221[0]), .Y(i_0_not_high_prior_arbiter1221) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1221), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1221[0]), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b1), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(_sv2v_jump_high_prior_arbiter1221[1]), .QN(nandres_high_prior_arbiter1221) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22212) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2221[0]), .Y(i_0_not_high_prior_arbiter22212) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22212), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2221[0]), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(_sv2v_jump_high_prior_arbiter2221[1]), .QN(nandres_high_prior_arbiter22212) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter221[0]), .B(valid_from_im_output_module2[7:4][0]), .Y(mask_req_rr_arbiter221[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter221[1]), .B(valid_from_im_output_module2[7:4][1]), .Y(mask_req_rr_arbiter221[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter221[0]), .Y(next_mask_rr_arbiter221[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter221[1]), .Y(next_mask_rr_arbiter221[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter221[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter221) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter221[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter221) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter221[0]), .IN2(raw_grant_rr_arbiter221[0]), .S(xnor0res_rr_arbiter221), .Q(grant_im_output_module2[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter221[1]), .IN2(raw_grant_rr_arbiter221[1]), .S(xnor1res_rr_arbiter221), .Q(grant_im_output_module2[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter221[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter221[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter221[1]), .B(1'b0), .Y(firstif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter221), .B(grant_im_output_module2[7:4][i_rr_arbiter221[0]]), .Y(secondif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[1]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter221[0]), .Q(j_rr_arbiter221[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter221), .B(j_rr_arbiter221[0]), .Y(thirdif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter221[j_rr_arbiter221[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter221), .Q(next_mask_rr_arbiter221[j_rr_arbiter221[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b1), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(_sv2v_jump_rr_rr_arbiter221[1]), .QN(fourthif_rr_arbiter221) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter221) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter221) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter221[0]), .IN2(next_mask_rr_arbiter221[0]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter221[1]), .IN2(next_mask_rr_arbiter221[1]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter222211), .IN2(1'sb1), .S(arst_value_rr_arbiter221), .Q(mask_ff_rr_arbiter221[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter1222[0]), .Y(i_0_not_high_prior_arbiter1222) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1222), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1222[0]), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b1), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(_sv2v_jump_high_prior_arbiter1222[1]), .QN(nandres_high_prior_arbiter1222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2222) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter2222[0]), .Y(i_0_not_high_prior_arbiter2222) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2222), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2222[0]), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(_sv2v_jump_high_prior_arbiter2222[1]), .QN(nandres_high_prior_arbiter2222) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter222[0]), .B(valid_from_im_output_module2[11:8][0]), .Y(mask_req_rr_arbiter222[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter222[1]), .B(valid_from_im_output_module2[11:8][1]), .Y(mask_req_rr_arbiter222[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter222[0]), .Y(next_mask_rr_arbiter222[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter222[1]), .Y(next_mask_rr_arbiter222[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter222[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter222) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter222[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter222) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter222[0]), .IN2(raw_grant_rr_arbiter222[0]), .S(xnor0res_rr_arbiter222), .Q(grant_im_output_module2[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter222[1]), .IN2(raw_grant_rr_arbiter222[1]), .S(xnor1res_rr_arbiter222), .Q(grant_im_output_module2[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter222[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter222[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter222[1]), .B(1'b0), .Y(firstif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter222), .B(grant_im_output_module2[11:8][i_rr_arbiter222[0]]), .Y(secondif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[1]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter222[0]), .Q(j_rr_arbiter222[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter222), .B(j_rr_arbiter222[0]), .Y(thirdif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter222[j_rr_arbiter222[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter222), .Q(next_mask_rr_arbiter222[j_rr_arbiter222[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b1), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(_sv2v_jump_rr_rr_arbiter222[1]), .QN(fourthif_rr_arbiter222) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter222) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter222) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter222[0]), .IN2(next_mask_rr_arbiter222[0]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter222[1]), .IN2(next_mask_rr_arbiter222[1]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter222222), .IN2(1'sb1), .S(arst_value_rr_arbiter222), .Q(mask_ff_rr_arbiter222[0]));


    XNOR2X1 U222 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37]), .IN2(vc_channel_output_module2[1]), .QN(xnor1resu1_output_module2) );
    XNOR2X1 U223 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37-1]), .IN2(vc_channel_output_module2[0]), .QN(xnor2resu1_output_module2) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module2), .IN2(xnor2resu1_output_module2), .Q(and1resu1_output_module2) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]), .IN2(1'b1), .S(and1resu1_output_module2), .Q(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .Q(xor1resu1_output_module2) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module2_1[0]), .IN2(_sv2v_jump_output_module2[0]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module2_1[1]), .IN2(_sv2v_jump_output_module2[1]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[vc_channel_output_module2[1:0]*4+in_mod_output_module2[1:0]]), .Q(and2resu1_output_module2) );

    MUX21X1 U3(.IN1(head_flit_output_module2[3]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+3]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[3]));
    MUX21X1 U4(.IN1(head_flit_output_module2[4]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+4]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[4]));
    MUX21X1 U5(.IN1(head_flit_output_module2[5]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+5]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[5]));
    MUX21X1 U6(.IN1(head_flit_output_module2[6]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+6]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[6]));
    MUX21X1 U7(.IN1(head_flit_output_module2[7]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+7]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[7]));
    MUX21X1 U8(.IN1(head_flit_output_module2[8]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+8]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[8]));
    MUX21X1 U9(.IN1(head_flit_output_module2[9]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+9]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[9]));
    MUX21X1 U10(.IN1(head_flit_output_module2[10]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+10]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[10]));
    MUX21X1 U11(.IN1(head_flit_output_module2[11]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+11]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[11]));
    MUX21X1 U12(.IN1(head_flit_output_module2[12]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+12]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[12]));
    MUX21X1 U13(.IN1(head_flit_output_module2[13]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+13]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[13]));
    MUX21X1 U14(.IN1(head_flit_output_module2[14]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+14]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[14]));
    MUX21X1 U15(.IN1(head_flit_output_module2[15]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+15]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[15]));
    MUX21X1 U16(.IN1(head_flit_output_module2[16]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+16]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[16]));
    MUX21X1 U17(.IN1(head_flit_output_module2[17]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+17]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[17]));
    MUX21X1 U18(.IN1(head_flit_output_module2[18]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+18]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[18]));
    MUX21X1 U19(.IN1(head_flit_output_module2[19]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+19]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[19]));
    MUX21X1 U20(.IN1(head_flit_output_module2[20]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+20]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[20]));
    MUX21X1 U21(.IN1(head_flit_output_module2[21]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+21]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[21]));
    MUX21X1 U22(.IN1(head_flit_output_module2[22]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+22]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[22]));
    MUX21X1 U23(.IN1(head_flit_output_module2[23]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+23]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[23]));
    MUX21X1 U24(.IN1(head_flit_output_module2[24]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+24]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[24]));
    MUX21X1 U25(.IN1(head_flit_output_module2[25]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+25]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[25]));
    MUX21X1 U26(.IN1(head_flit_output_module2[26]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+26]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[26]));
    MUX21X1 U27(.IN1(head_flit_output_module2[27]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+27]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[27]));
    MUX21X1 U28(.IN1(head_flit_output_module2[28]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+28]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[28]));
    MUX21X1 U29(.IN1(head_flit_output_module2[29]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+29]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[29]));
    MUX21X1 U30(.IN1(head_flit_output_module2[30]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+30]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[30]));
    MUX21X1 U31(.IN1(head_flit_output_module2[31]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+31]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[31]));
    MUX21X1 U32(.IN1(head_flit_output_module2[32]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+32]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[32]));
    MUX21X1 U33(.IN1(head_flit_output_module2[33]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+33]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[33]));
    MUX21X1 U34(.IN1(head_flit_output_module2[34]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+34]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[34]));
    MUX21X1 U35(.IN1(head_flit_output_module2[35]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+35]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[35]));
    MUX21X1 U36(.IN1(head_flit_output_module2[36]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+36]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[36]));

    INVX1 U041 ( .A(head_flit_output_module2[32]), .Y(head_flit_output_module2_32_not_output_module2) );
    AND2X1 U1218 ( .IN1(head_flit_output_module2_32_not_output_module2), .IN2(head_flit_output_module2[33]), .Q(and3resu1_output_module2) );
    NOR4X1 U175821 (.IN1(head_flit_output_module2[29]), .IN2(head_flit_output_module2[28]), .IN3(head_flit_output_module2[27]), .IN4(head_flit_output_module2[26]), .Q(nor23resu1_output_module2) );
    NOR4X1 U175831 (.IN1(head_flit_output_module2[25]), .IN2(head_flit_output_module2[24]), .IN3(head_flit_output_module2[23]), .IN4(head_flit_output_module2[22]), .Q(nor23resu2_output_module2) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module2), .IN2(nor23resu2_output_module2), .Q(and4resu1_output_module2) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module2[33]), .IN2(head_flit_output_module2[32]), .Q(nor23resu3_output_module2) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module2), .IN2(and4resu1_output_module2), .Q(and5resu1_output_module2) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module2), .IN2(nor23resu3_output_module2), .Q(or12resu12_output_module2) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[3:2][0]), .IN2(or12resu12_output_module2), .Q(and6resu1_output_module2) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]), .IN2(and6resu1_output_module2), .S(and2resu1_output_module2) ,.Q(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module2[0]),.B(_sv2v_jump_output_module2[1]),.Y(nand1resu_output_module2));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(_sv2v_jump_output_module2_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module2[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module2[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[i_output_module2[1:0] * 4+:4]), .Q(and8resu1_output_module2) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module2[0]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module2[1]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[1]);
    MUX21X1 U3631(.IN1(req_out_output_module2), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(req_out_output_module2);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2[1]), .Q(norfinresu1_output_module2) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module2), .IN2(req_out_output_module2), .Q(and9resu1_output_module2) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module2), .IN2(grant_im_output_module2[(vc_ch_act_out_output_module2 * 4) + i_output_module2[1:0]]), .Q(and10resu1_output_module2) );    

    MUX21X1 U3(.IN1(ext_req_v_o[110:74][3]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+3]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[110:74][4]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+4]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[110:74][5]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+5]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[110:74][6]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+6]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[110:74][7]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+7]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[110:74][8]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+8]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[110:74][9]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+9]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[110:74][10]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+10]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[110:74][11]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+11]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[110:74][12]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+12]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[110:74][13]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+13]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[110:74][14]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+14]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[110:74][15]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+15]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[110:74][16]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+16]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[110:74][17]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+17]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[110:74][18]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+18]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[110:74][19]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+19]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[110:74][20]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+20]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[110:74][21]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+21]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[110:74][22]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+22]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[110:74][23]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+23]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[110:74][24]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+24]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[110:74][25]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+25]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[110:74][26]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+26]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[110:74][27]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+27]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[110:74][28]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+28]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[110:74][29]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+29]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[110:74][30]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+30]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[110:74][31]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+31]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[110:74][32]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+32]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[110:74][33]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+33]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[110:74][34]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+34]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[110:74][35]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+35]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[110:74][36]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+36]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[110:74][0]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[110:74][1]), .IN2(vc_ch_act_out_output_module2[0]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[110:74][2]), .IN2(vc_ch_act_out_output_module2[1]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and11resu1_output_module2) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);   










    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter13) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter13[0]), .Y(i_0_not_high_prior_arbiter13) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter13), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter13[0]), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b1), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(_sv2v_jump_high_prior_arbiter13[1]), .QN(nandres_high_prior_arbiter13) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter23) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter23[0]), .Y(i_0_not_high_prior_arbiter23) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter23), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter23[0]), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(_sv2v_jump_high_prior_arbiter23[1]), .QN(nandres_high_prior_arbiter23) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter3[0]), .B(valid_from_im_output_module3[3:0][0]), .Y(mask_req_rr_arbiter3[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter3[1]), .B(valid_from_im_output_module3[3:0][1]), .Y(mask_req_rr_arbiter3[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter3[0]), .Y(next_mask_rr_arbiter3[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter3[1]), .Y(next_mask_rr_arbiter3[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter3[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter3) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter3[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter3) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter3[0]), .IN2(raw_grant_rr_arbiter3[0]), .S(xnor0res_rr_arbiter3), .Q(grant_im_output_module3[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter3[1]), .IN2(raw_grant_rr_arbiter3[1]), .S(xnor1res_rr_arbiter3), .Q(grant_im_output_module3[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter3[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter3[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter3[1]), .B(1'b0), .Y(firstif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter3), .B(grant_im_output_module3[3:0][i_rr_arbiter3[0]]), .Y(secondif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[1]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter3[0]), .Q(j_rr_arbiter3[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter3), .B(j_rr_arbiter3[0]), .Y(thirdif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter3[j_rr_arbiter3[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter3), .Q(next_mask_rr_arbiter3[j_rr_arbiter3[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b1), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(_sv2v_jump_rr_rr_arbiter3[1]), .QN(fourthif_rr_arbiter3) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter3) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter3) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter3[0]), .IN2(next_mask_rr_arbiter3[0]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter3[1]), .IN2(next_mask_rr_arbiter3[1]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter33), .IN2(1'sb1), .S(arst_value_rr_arbiter3), .Q(mask_ff_rr_arbiter3[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter131) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter131[0]), .Y(i_0_not_high_prior_arbiter131) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter131), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter131[0]), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b1), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(_sv2v_jump_high_prior_arbiter131[1]), .QN(nandres_high_prior_arbiter131) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2313) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter231[0]), .Y(i_0_not_high_prior_arbiter2313) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2313), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter231[0]), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(_sv2v_jump_high_prior_arbiter231[1]), .QN(nandres_high_prior_arbiter2313) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter31[0]), .B(valid_from_im_output_module3[7:4][0]), .Y(mask_req_rr_arbiter31[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter31[1]), .B(valid_from_im_output_module3[7:4][1]), .Y(mask_req_rr_arbiter31[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter31[0]), .Y(next_mask_rr_arbiter31[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter31[1]), .Y(next_mask_rr_arbiter31[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter31[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter31) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter31[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter31) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter31[0]), .IN2(raw_grant_rr_arbiter31[0]), .S(xnor0res_rr_arbiter31), .Q(grant_im_output_module3[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter31[1]), .IN2(raw_grant_rr_arbiter31[1]), .S(xnor1res_rr_arbiter31), .Q(grant_im_output_module3[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter31[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter31[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter31[1]), .B(1'b0), .Y(firstif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter31), .B(grant_im_output_module3[7:4][i_rr_arbiter31[0]]), .Y(secondif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[1]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter31[0]), .Q(j_rr_arbiter31[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter31), .B(j_rr_arbiter31[0]), .Y(thirdif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter31[j_rr_arbiter31[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter31), .Q(next_mask_rr_arbiter31[j_rr_arbiter31[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b1), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(_sv2v_jump_rr_rr_arbiter31[1]), .QN(fourthif_rr_arbiter31) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter31) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter31) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter31[0]), .IN2(next_mask_rr_arbiter31[0]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter31[1]), .IN2(next_mask_rr_arbiter31[1]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter3311), .IN2(1'sb1), .S(arst_value_rr_arbiter31), .Q(mask_ff_rr_arbiter31[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter132) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter132[0]), .Y(i_0_not_high_prior_arbiter132) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter132), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter132[0]), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b1), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(_sv2v_jump_high_prior_arbiter132[1]), .QN(nandres_high_prior_arbiter132) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter232) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter232[0]), .Y(i_0_not_high_prior_arbiter232) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter232), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter232[0]), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(_sv2v_jump_high_prior_arbiter232[1]), .QN(nandres_high_prior_arbiter232) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter32[0]), .B(valid_from_im_output_module3[11:8][0]), .Y(mask_req_rr_arbiter32[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter32[1]), .B(valid_from_im_output_module3[11:8][1]), .Y(mask_req_rr_arbiter32[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter32[0]), .Y(next_mask_rr_arbiter32[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter32[1]), .Y(next_mask_rr_arbiter32[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter32[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter32) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter32[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter32) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter32[0]), .IN2(raw_grant_rr_arbiter32[0]), .S(xnor0res_rr_arbiter32), .Q(grant_im_output_module3[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter32[1]), .IN2(raw_grant_rr_arbiter32[1]), .S(xnor1res_rr_arbiter32), .Q(grant_im_output_module3[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter32[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter32[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter32[1]), .B(1'b0), .Y(firstif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter32), .B(grant_im_output_module3[11:8][i_rr_arbiter32[0]]), .Y(secondif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[1]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter32[0]), .Q(j_rr_arbiter32[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter32), .B(j_rr_arbiter32[0]), .Y(thirdif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter32[j_rr_arbiter32[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter32), .Q(next_mask_rr_arbiter32[j_rr_arbiter32[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b1), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(_sv2v_jump_rr_rr_arbiter32[1]), .QN(fourthif_rr_arbiter32) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter32) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter32) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter32[0]), .IN2(next_mask_rr_arbiter32[0]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter32[1]), .IN2(next_mask_rr_arbiter32[1]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter3322), .IN2(1'sb1), .S(arst_value_rr_arbiter32), .Q(mask_ff_rr_arbiter32[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37]), .IN2(vc_channel_output_module3[1]), .QN(xnor1resu1_output_module3) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37-1]), .IN2(vc_channel_output_module3[0]), .QN(xnor2resu1_output_module3) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module3), .IN2(xnor2resu1_output_module3), .Q(and1resu1_output_module3) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]), .IN2(1'b1), .S(and1resu1_output_module3), .Q(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .Q(xor1resu1_output_module3) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module3_1[0]), .IN2(_sv2v_jump_output_module3[0]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module3_1[1]), .IN2(_sv2v_jump_output_module3[1]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[vc_channel_output_module3[1:0]*4+in_mod_output_module3[1:0]]), .Q(and2resu1_output_module3) );

    MUX21X1 U3(.IN1(head_flit_output_module3[3]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+3]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[3]));
    MUX21X1 U4(.IN1(head_flit_output_module3[4]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+4]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[4]));
    MUX21X1 U5(.IN1(head_flit_output_module3[5]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+5]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[5]));
    MUX21X1 U6(.IN1(head_flit_output_module3[6]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+6]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[6]));
    MUX21X1 U7(.IN1(head_flit_output_module3[7]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+7]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[7]));
    MUX21X1 U8(.IN1(head_flit_output_module3[8]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+8]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[8]));
    MUX21X1 U9(.IN1(head_flit_output_module3[9]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+9]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[9]));
    MUX21X1 U10(.IN1(head_flit_output_module3[10]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+10]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[10]));
    MUX21X1 U11(.IN1(head_flit_output_module3[11]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+11]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[11]));
    MUX21X1 U12(.IN1(head_flit_output_module3[12]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+12]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[12]));
    MUX21X1 U13(.IN1(head_flit_output_module3[13]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+13]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[13]));
    MUX21X1 U14(.IN1(head_flit_output_module3[14]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+14]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[14]));
    MUX21X1 U15(.IN1(head_flit_output_module3[15]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+15]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[15]));
    MUX21X1 U16(.IN1(head_flit_output_module3[16]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+16]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[16]));
    MUX21X1 U17(.IN1(head_flit_output_module3[17]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+17]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[17]));
    MUX21X1 U18(.IN1(head_flit_output_module3[18]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+18]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[18]));
    MUX21X1 U19(.IN1(head_flit_output_module3[19]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+19]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[19]));
    MUX21X1 U20(.IN1(head_flit_output_module3[20]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+20]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[20]));
    MUX21X1 U21(.IN1(head_flit_output_module3[21]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+21]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[21]));
    MUX21X1 U22(.IN1(head_flit_output_module3[22]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+22]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[22]));
    MUX21X1 U23(.IN1(head_flit_output_module3[23]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+23]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[23]));
    MUX21X1 U24(.IN1(head_flit_output_module3[24]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+24]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[24]));
    MUX21X1 U25(.IN1(head_flit_output_module3[25]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+25]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[25]));
    MUX21X1 U26(.IN1(head_flit_output_module3[26]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+26]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[26]));
    MUX21X1 U27(.IN1(head_flit_output_module3[27]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+27]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[27]));
    MUX21X1 U28(.IN1(head_flit_output_module3[28]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+28]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[28]));
    MUX21X1 U29(.IN1(head_flit_output_module3[29]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+29]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[29]));
    MUX21X1 U30(.IN1(head_flit_output_module3[30]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+30]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[30]));
    MUX21X1 U31(.IN1(head_flit_output_module3[31]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+31]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[31]));
    MUX21X1 U32(.IN1(head_flit_output_module3[32]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+32]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[32]));
    MUX21X1 U33(.IN1(head_flit_output_module3[33]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+33]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[33]));
    MUX21X1 U34(.IN1(head_flit_output_module3[34]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+34]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[34]));
    MUX21X1 U35(.IN1(head_flit_output_module3[35]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+35]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[35]));
    MUX21X1 U36(.IN1(head_flit_output_module3[36]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+36]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[36]));

    INVX1 U041 ( .A(head_flit_output_module3[32]), .Y(head_flit_output_module3_32_not_output_module3) );
    AND2X1 U1218 ( .IN1(head_flit_output_module3_32_not_output_module3), .IN2(head_flit_output_module3[33]), .Q(and3resu1_output_module3) );
    NOR4X1 U175821 (.IN1(head_flit_output_module3[29]), .IN2(head_flit_output_module3[28]), .IN3(head_flit_output_module3[27]), .IN4(head_flit_output_module3[26]), .Q(nor23resu1_output_module3) );
    NOR4X1 U175831 (.IN1(head_flit_output_module3[25]), .IN2(head_flit_output_module3[24]), .IN3(head_flit_output_module3[23]), .IN4(head_flit_output_module3[22]), .Q(nor23resu2_output_module3) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module3), .IN2(nor23resu2_output_module3), .Q(and4resu1_output_module3) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module3[33]), .IN2(head_flit_output_module3[32]), .Q(nor23resu3_output_module3) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module3), .IN2(and4resu1_output_module3), .Q(and5resu1_output_module3) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module3), .IN2(nor23resu3_output_module3), .Q(or12resu12_output_module3) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[4:3][0]), .IN2(or12resu12_output_module3), .Q(and6resu1_output_module3) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]), .IN2(and6resu1_output_module3), .S(and2resu1_output_module3) ,.Q(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module3[0]),.B(_sv2v_jump_output_module3[1]),.Y(nand1resu_output_module3));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(_sv2v_jump_output_module3_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module3[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module3[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[i_output_module3[1:0] * 4+:4]), .Q(and8resu1_output_module3) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module3[0]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module3[1]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[1]);
    MUX21X1 U3631(.IN1(req_out_output_module3), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(req_out_output_module3);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3[1]), .Q(norfinresu1_output_module3) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module3), .IN2(req_out_output_module3), .Q(and9resu1_output_module3) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module3), .IN2(grant_im_output_module3[(vc_ch_act_out_output_module3 * 4) + i_output_module3[1:0]]), .Q(and10resu1_output_module3) );    

    MUX21X1 U3(.IN1(ext_req_v_o[147:111][3]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+3]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[147:111][4]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+4]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[147:111][5]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+5]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[147:111][6]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+6]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[147:111][7]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+7]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[147:111][8]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+8]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[147:111][9]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+9]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[147:111][10]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+10]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[147:111][11]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+11]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[147:111][12]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+12]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[147:111][13]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+13]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[147:111][14]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+14]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[147:111][15]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+15]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[147:111][16]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+16]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[147:111][17]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+17]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[147:111][18]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+18]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[147:111][19]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+19]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[147:111][20]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+20]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[147:111][21]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+21]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[147:111][22]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+22]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[147:111][23]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+23]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[147:111][24]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+24]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[147:111][25]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+25]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[147:111][26]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+26]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[147:111][27]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+27]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[147:111][28]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+28]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[147:111][29]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+29]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[147:111][30]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+30]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[147:111][31]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+31]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[147:111][32]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+32]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[147:111][33]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+33]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[147:111][34]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+34]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[147:111][35]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+35]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[147:111][36]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+36]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[147:111][0]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[147:111][1]), .IN2(vc_ch_act_out_output_module3[0]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[147:111][2]), .IN2(vc_ch_act_out_output_module3[1]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and11resu1_output_module3) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    







    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter14) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter14[0]), .Y(i_0_not_high_prior_arbiter14) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter14), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter14[0]), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b1), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(_sv2v_jump_high_prior_arbiter14[1]), .QN(nandres_high_prior_arbiter14) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter24) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter24[0]), .Y(i_0_not_high_prior_arbiter24) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter24), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter24[0]), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(_sv2v_jump_high_prior_arbiter24[1]), .QN(nandres_high_prior_arbiter24) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter4[0]), .B(valid_from_im_output_module4[3:0][0]), .Y(mask_req_rr_arbiter4[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter4[1]), .B(valid_from_im_output_module4[3:0][1]), .Y(mask_req_rr_arbiter4[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter4[0]), .Y(next_mask_rr_arbiter4[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter4[1]), .Y(next_mask_rr_arbiter4[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter4[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter4) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter4[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter4) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter4[0]), .IN2(raw_grant_rr_arbiter4[0]), .S(xnor0res_rr_arbiter4), .Q(grant_im_output_module4[3:0][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter4[1]), .IN2(raw_grant_rr_arbiter4[1]), .S(xnor1res_rr_arbiter4), .Q(grant_im_output_module4[3:0][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter4[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter4[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter4[1]), .B(1'b0), .Y(firstif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter4), .B(grant_im_output_module4[3:0][i_rr_arbiter4[0]]), .Y(secondif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[1]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter4[0]), .Q(j_rr_arbiter4[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter4), .B(j_rr_arbiter4[0]), .Y(thirdif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter4[j_rr_arbiter4[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter4), .Q(next_mask_rr_arbiter4[j_rr_arbiter4[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b1), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(_sv2v_jump_rr_rr_arbiter4[1]), .QN(fourthif_rr_arbiter4) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter4) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter4) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter4[0]), .IN2(next_mask_rr_arbiter4[0]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter4[1]), .IN2(next_mask_rr_arbiter4[1]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter44), .IN2(1'sb1), .S(arst_value_rr_arbiter4), .Q(mask_ff_rr_arbiter4[0]));



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter141) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter141[0]), .Y(i_0_not_high_prior_arbiter141) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter141), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter141[0]), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b1), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(_sv2v_jump_high_prior_arbiter141[1]), .QN(nandres_high_prior_arbiter141) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2414) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter241[0]), .Y(i_0_not_high_prior_arbiter2414) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2414), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter241[0]), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(_sv2v_jump_high_prior_arbiter241[1]), .QN(nandres_high_prior_arbiter2414) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter41[0]), .B(valid_from_im_output_module4[7:4][0]), .Y(mask_req_rr_arbiter41[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter41[1]), .B(valid_from_im_output_module4[7:4][1]), .Y(mask_req_rr_arbiter41[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter41[0]), .Y(next_mask_rr_arbiter41[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter41[1]), .Y(next_mask_rr_arbiter41[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter41[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter41) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter41[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter41) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter41[0]), .IN2(raw_grant_rr_arbiter41[0]), .S(xnor0res_rr_arbiter41), .Q(grant_im_output_module4[7:4][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter41[1]), .IN2(raw_grant_rr_arbiter41[1]), .S(xnor1res_rr_arbiter41), .Q(grant_im_output_module4[7:4][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter41[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter41[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter41[1]), .B(1'b0), .Y(firstif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter41), .B(grant_im_output_module4[7:4][i_rr_arbiter41[0]]), .Y(secondif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[1]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter41[0]), .Q(j_rr_arbiter41[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter41), .B(j_rr_arbiter41[0]), .Y(thirdif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter41[j_rr_arbiter41[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter41), .Q(next_mask_rr_arbiter41[j_rr_arbiter41[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b1), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(_sv2v_jump_rr_rr_arbiter41[1]), .QN(fourthif_rr_arbiter41) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter41) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter41) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter41[0]), .IN2(next_mask_rr_arbiter41[0]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter41[1]), .IN2(next_mask_rr_arbiter41[1]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter4411), .IN2(1'sb1), .S(arst_value_rr_arbiter41), .Q(mask_ff_rr_arbiter41[0]));





    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter142) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter142[0]), .Y(i_0_not_high_prior_arbiter142) );
    MUX21X1 U09 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter142), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[0]);
    MUX21X1 U10 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter142[0]), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b1), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(_sv2v_jump_high_prior_arbiter142[1]), .QN(nandres_high_prior_arbiter142) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );



    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[1]) );
    BUFX1 U02 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U03 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    XNOR2X1 U05 ( .IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter242) );
    MUX21X1 U06 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U07 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    INVX1 U08 ( .A(i_high_prior_arbiter242[0]), .Y(i_0_not_high_prior_arbiter242) );
    MUX21X1 U09 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter242), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[0]);
    MUX21X1 U10 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter242[0]), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[1]);
    MUX21X1 U11 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U12 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    NAND2X1 U13 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(_sv2v_jump_high_prior_arbiter242[1]), .QN(nandres_high_prior_arbiter242) );
    MUX21X1 U14 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U15 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    HADDX1 U00021 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U00022 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U00021 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    

    BUFX1 U00 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[0]) );
    BUFX1 U01 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[1]) );
    AND2X1 U02 ( .A(mask_ff_rr_arbiter42[0]), .B(valid_from_im_output_module4[11:8][0]), .Y(mask_req_rr_arbiter42[0]) );
    AND2X1 U03 ( .A(mask_ff_rr_arbiter42[1]), .B(valid_from_im_output_module4[11:8][1]), .Y(mask_req_rr_arbiter42[1]) );
    BUFX1 U04 ( .A(mask_ff_rr_arbiter42[0]), .Y(next_mask_rr_arbiter42[0]) );
    BUFX1 U05 ( .A(mask_ff_rr_arbiter42[1]), .Y(next_mask_rr_arbiter42[1]) );
    XNOR2X1 U06 ( .IN1(mask_req_rr_arbiter42[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter42) );
    XNOR2X1 U07 ( .IN1(mask_req_rr_arbiter42[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter42) );
    MUX21X1 U08 (.IN1(masked_grant_rr_arbiter42[0]), .IN2(raw_grant_rr_arbiter42[0]), .S(xnor0res_rr_arbiter42), .Q(grant_im_output_module4[11:8][0]));
    MUX21X1 U09 (.IN1(masked_grant_rr_arbiter42[1]), .IN2(raw_grant_rr_arbiter42[1]), .S(xnor1res_rr_arbiter42), .Q(grant_im_output_module4[11:8][1]));

    BUFX1 U00 ( .A(1'b0), .Y(i_rr_arbiter42[1]) );
    MUX21X1 U09 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter42[0]));

    AND2X1 U02 ( .A(_sv2v_jump_rr_rr_arbiter42[1]), .B(1'b0), .Y(firstif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    AND2X1 U02 ( .A(firstif_rr_arbiter42), .B(grant_im_output_module4[11:8][i_rr_arbiter42[0]]), .Y(secondif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[1]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[1]));
    MUX21X1 U09 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter42[0]), .Q(j_rr_arbiter42[0]));
    AND2X1 U02 ( .A(secondif_rr_arbiter42), .B(j_rr_arbiter42[0]), .Y(thirdif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(next_mask_rr_arbiter42[j_rr_arbiter42[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter42), .Q(next_mask_rr_arbiter42[j_rr_arbiter42[0]]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b1), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    NAND2X1 U213 ( .IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(_sv2v_jump_rr_rr_arbiter42[1]), .QN(fourthif_rr_arbiter42) );
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    MUX21X1 U09 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    DFFX2 U30 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter42) );
    DFFX2 U31 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter42) );
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter42[0]), .IN2(next_mask_rr_arbiter42[0]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[0]));
    MUX21X1 U09 (.IN1(mask_ff_rr_arbiter42[1]), .IN2(next_mask_rr_arbiter42[1]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[1]));
    MUX21X1 U09 (.IN1(temp_mask_ff_rr_arbiter4422), .IN2(1'sb1), .S(arst_value_rr_arbiter42), .Q(mask_ff_rr_arbiter42[0]));


    XNOR2X1 U222 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37]), .IN2(vc_channel_output_module4[1]), .QN(xnor1resu1_output_module4) );
    XNOR2X1 U223 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37-1]), .IN2(vc_channel_output_module4[0]), .QN(xnor2resu1_output_module4) );
    AND2X1 U128 ( .IN1(xnor1resu1_output_module4), .IN2(xnor2resu1_output_module4), .Q(and1resu1_output_module4) );
    MUX21X1 U0009 (.IN1(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]), .IN2(1'b1), .S(and1resu1_output_module4), .Q(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]);
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );  
    HADDX1 U00023 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00022 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) ); 
    XOR2X1 U02221 ( .IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .Q(xor1resu1_output_module4) );
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[1]));
    MUX21X1 U00171 (.IN1(_sv2v_jump_output_module4_1[0]), .IN2(_sv2v_jump_output_module4[0]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[0]));
    MUX21X1 U00181 (.IN1(_sv2v_jump_output_module4_1[1]), .IN2(_sv2v_jump_output_module4[1]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[1]));
    AND2X1 U1218 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[vc_channel_output_module4[1:0]*4+in_mod_output_module4[1:0]]), .Q(and2resu1_output_module4) );

    MUX21X1 U3(.IN1(head_flit_output_module4[3]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+3]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[3]));
    MUX21X1 U4(.IN1(head_flit_output_module4[4]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+4]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[4]));
    MUX21X1 U5(.IN1(head_flit_output_module4[5]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+5]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[5]));
    MUX21X1 U6(.IN1(head_flit_output_module4[6]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+6]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[6]));
    MUX21X1 U7(.IN1(head_flit_output_module4[7]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+7]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[7]));
    MUX21X1 U8(.IN1(head_flit_output_module4[8]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+8]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[8]));
    MUX21X1 U9(.IN1(head_flit_output_module4[9]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+9]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[9]));
    MUX21X1 U10(.IN1(head_flit_output_module4[10]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+10]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[10]));
    MUX21X1 U11(.IN1(head_flit_output_module4[11]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+11]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[11]));
    MUX21X1 U12(.IN1(head_flit_output_module4[12]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+12]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[12]));
    MUX21X1 U13(.IN1(head_flit_output_module4[13]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+13]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[13]));
    MUX21X1 U14(.IN1(head_flit_output_module4[14]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+14]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[14]));
    MUX21X1 U15(.IN1(head_flit_output_module4[15]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+15]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[15]));
    MUX21X1 U16(.IN1(head_flit_output_module4[16]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+16]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[16]));
    MUX21X1 U17(.IN1(head_flit_output_module4[17]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+17]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[17]));
    MUX21X1 U18(.IN1(head_flit_output_module4[18]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+18]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[18]));
    MUX21X1 U19(.IN1(head_flit_output_module4[19]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+19]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[19]));
    MUX21X1 U20(.IN1(head_flit_output_module4[20]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+20]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[20]));
    MUX21X1 U21(.IN1(head_flit_output_module4[21]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+21]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[21]));
    MUX21X1 U22(.IN1(head_flit_output_module4[22]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+22]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[22]));
    MUX21X1 U23(.IN1(head_flit_output_module4[23]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+23]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[23]));
    MUX21X1 U24(.IN1(head_flit_output_module4[24]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+24]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[24]));
    MUX21X1 U25(.IN1(head_flit_output_module4[25]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+25]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[25]));
    MUX21X1 U26(.IN1(head_flit_output_module4[26]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+26]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[26]));
    MUX21X1 U27(.IN1(head_flit_output_module4[27]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+27]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[27]));
    MUX21X1 U28(.IN1(head_flit_output_module4[28]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+28]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[28]));
    MUX21X1 U29(.IN1(head_flit_output_module4[29]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+29]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[29]));
    MUX21X1 U30(.IN1(head_flit_output_module4[30]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+30]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[30]));
    MUX21X1 U31(.IN1(head_flit_output_module4[31]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+31]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[31]));
    MUX21X1 U32(.IN1(head_flit_output_module4[32]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+32]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[32]));
    MUX21X1 U33(.IN1(head_flit_output_module4[33]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+33]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[33]));
    MUX21X1 U34(.IN1(head_flit_output_module4[34]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+34]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[34]));
    MUX21X1 U35(.IN1(head_flit_output_module4[35]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+35]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[35]));
    MUX21X1 U36(.IN1(head_flit_output_module4[36]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+36]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[36]));

    INVX1 U041 ( .A(head_flit_output_module4[32]), .Y(head_flit_output_module4_32_not_output_module4) );
    AND2X1 U1218 ( .IN1(head_flit_output_module4_32_not_output_module4), .IN2(head_flit_output_module4[33]), .Q(and3resu1_output_module4) );
    NOR4X1 U175821 (.IN1(head_flit_output_module4[29]), .IN2(head_flit_output_module4[28]), .IN3(head_flit_output_module4[27]), .IN4(head_flit_output_module4[26]), .Q(nor23resu1_output_module4) );
    NOR4X1 U175831 (.IN1(head_flit_output_module4[25]), .IN2(head_flit_output_module4[24]), .IN3(head_flit_output_module4[23]), .IN4(head_flit_output_module4[22]), .Q(nor23resu2_output_module4) );
    AND2X1 U12183 ( .IN1(nor23resu1_output_module4), .IN2(nor23resu2_output_module4), .Q(and4resu1_output_module4) );
    NOR2X1 U1758211 (.IN1(head_flit_output_module4[33]), .IN2(head_flit_output_module4[32]), .Q(nor23resu3_output_module4) );
    AND2X1 U12183 ( .IN1(nor23resu3_output_module4), .IN2(and4resu1_output_module4), .Q(and5resu1_output_module4) );    
    OR2X1 U17582121 (.IN1(and3resu1_output_module4), .IN2(nor23resu3_output_module4), .Q(or12resu12_output_module4) );
    AND2X1 U12183 ( .IN1(ext_resp_v_i[5:4][0]), .IN2(or12resu12_output_module4), .Q(and6resu1_output_module4) );    
    MUX21X1 U361(.IN1(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]), .IN2(and6resu1_output_module4), .S(and2resu1_output_module4) ,.Q(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    NAND2X1 U29311(.A(_sv2v_jump_output_module4[0]),.B(_sv2v_jump_output_module4[1]),.Y(nand1resu_output_module4));

    AND2X1 U12483 ( .IN1(xor1resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and7resu1) );    
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(_sv2v_jump_output_module4_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );



    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module4[0]));
    BUFX1 U4(.A(1'b0), .Y(_sv2v_jump_output_module4[1]));
    AND2X1 U12483 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[i_output_module4[1:0] * 4+:4]), .Q(and8resu1_output_module4) );    
    MUX21X1 U3621(.IN1(vc_ch_act_out_output_module4[0]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[0]);
    MUX21X1 U3631(.IN1(vc_ch_act_out_output_module4[1]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[1]);
    MUX21X1 U3631(.IN1(req_out_output_module4), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(req_out_output_module4);
    MUX21X1 U3621(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U3631(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U00021 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );

    NOR2X1 U1758211 (.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4[1]), .Q(norfinresu1_output_module4) );
    AND2X1 U124831 ( .IN1(norfinresu1_output_module4), .IN2(req_out_output_module4), .Q(and9resu1_output_module4) );    
    HADDX1 U00021 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    AND2X1 U124831 ( .IN1(and9resu1_output_module4), .IN2(grant_im_output_module4[(vc_ch_act_out_output_module4 * 4) + i_output_module4[1:0]]), .Q(and10resu1_output_module4) );    

    MUX21X1 U3(.IN1(ext_req_v_o[184:148][3]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+3]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][3]));
    MUX21X1 U4(.IN1(ext_req_v_o[184:148][4]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+4]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][4]));
    MUX21X1 U5(.IN1(ext_req_v_o[184:148][5]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+5]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][5]));
    MUX21X1 U6(.IN1(ext_req_v_o[184:148][6]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+6]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][6]));
    MUX21X1 U7(.IN1(ext_req_v_o[184:148][7]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+7]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][7]));
    MUX21X1 U8(.IN1(ext_req_v_o[184:148][8]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+8]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][8]));
    MUX21X1 U9(.IN1(ext_req_v_o[184:148][9]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+9]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][9]));
    MUX21X1 U10(.IN1(ext_req_v_o[184:148][10]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+10]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][10]));
    MUX21X1 U11(.IN1(ext_req_v_o[184:148][11]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+11]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][11]));
    MUX21X1 U12(.IN1(ext_req_v_o[184:148][12]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+12]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][12]));
    MUX21X1 U13(.IN1(ext_req_v_o[184:148][13]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+13]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][13]));
    MUX21X1 U14(.IN1(ext_req_v_o[184:148][14]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+14]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][14]));
    MUX21X1 U15(.IN1(ext_req_v_o[184:148][15]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+15]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][15]));
    MUX21X1 U16(.IN1(ext_req_v_o[184:148][16]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+16]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][16]));
    MUX21X1 U17(.IN1(ext_req_v_o[184:148][17]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+17]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][17]));
    MUX21X1 U18(.IN1(ext_req_v_o[184:148][18]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+18]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][18]));
    MUX21X1 U19(.IN1(ext_req_v_o[184:148][19]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+19]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][19]));
    MUX21X1 U20(.IN1(ext_req_v_o[184:148][20]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+20]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][20]));
    MUX21X1 U21(.IN1(ext_req_v_o[184:148][21]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+21]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][21]));
    MUX21X1 U22(.IN1(ext_req_v_o[184:148][22]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+22]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][22]));
    MUX21X1 U23(.IN1(ext_req_v_o[184:148][23]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+23]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][23]));
    MUX21X1 U24(.IN1(ext_req_v_o[184:148][24]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+24]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][24]));
    MUX21X1 U25(.IN1(ext_req_v_o[184:148][25]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+25]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][25]));
    MUX21X1 U26(.IN1(ext_req_v_o[184:148][26]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+26]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][26]));
    MUX21X1 U27(.IN1(ext_req_v_o[184:148][27]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+27]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][27]));
    MUX21X1 U28(.IN1(ext_req_v_o[184:148][28]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+28]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][28]));
    MUX21X1 U29(.IN1(ext_req_v_o[184:148][29]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+29]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][29]));
    MUX21X1 U30(.IN1(ext_req_v_o[184:148][30]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+30]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][30]));
    MUX21X1 U31(.IN1(ext_req_v_o[184:148][31]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+31]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][31]));
    MUX21X1 U32(.IN1(ext_req_v_o[184:148][32]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+32]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][32]));
    MUX21X1 U33(.IN1(ext_req_v_o[184:148][33]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+33]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][33]));
    MUX21X1 U34(.IN1(ext_req_v_o[184:148][34]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+34]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][34]));
    MUX21X1 U35(.IN1(ext_req_v_o[184:148][35]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+35]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][35]));
    MUX21X1 U36(.IN1(ext_req_v_o[184:148][36]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+36]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][36]));

    MUX21X1 U36221(.IN1(ext_req_v_o[184:148][0]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][0]);
    MUX21X1 U36221(.IN1(ext_req_v_o[184:148][1]), .IN2(vc_ch_act_out_output_module4[0]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][1]);
    MUX21X1 U36331(.IN1(ext_req_v_o[184:148][2]), .IN2(vc_ch_act_out_output_module4[1]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][2]);    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    

    AND2X1 U124831 ( .IN1(and9resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and11resu1_output_module4) );    
    MUX21X1 U36221(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U36331(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    



//router body
	BUFX1 U001 ( .A(north_recv_req), .Y(ext_req_v_i[0]) );
	BUFX1 U002 ( .A(north_recv_resp), .Y(ext_resp_v_o[0]) );
	BUFX1 U003 ( .A(xt_req_v_i[37]), .Y(south_recv_req) );
	BUFX1 U004 ( .A(south_recv_resp), .Y(ext_resp_v_o[1]) );
	BUFX1 U005 ( .A(ext_req_v_i[74]), .Y(west_recv_req) );
	BUFX1 U006 ( .A(west_recv_resp), .Y(ext_resp_v_o[2]) );
	BUFX1 U007 ( .A(ext_req_v_i[111]), .Y(east_recv_req) );
	BUFX1 U008 ( .A(east_recv_resp), .Y(ext_resp_v_o[3]) );
	BUFX1 U009 ( .A(north_send_req), .Y(ext_req_v_o[0]) );
	BUFX1 U010 ( .A(ext_resp_v_i[0]), .Y(north_send_resp) );
	BUFX1 U011 ( .A(south_send_req), .Y(ext_req_v_o[37]) );
	BUFX1 U012 ( .A(ext_resp_v_i[1]), .Y(south_send_resp) );
	BUFX1 U013 ( .A(west_send_req), .Y(ext_req_v_o[74]) );
	BUFX1 U014 ( .A(ext_resp_v_i[2]), .Y(west_send_resp) );
	BUFX1 U015 ( .A(east_send_req), .Y(ext_req_v_o[111]) );
	BUFX1 U016 ( .A(ext_resp_v_i[3]), .Y(east_send_resp) );
	BUFX1 U017 ( .A(local_recv_resp), .Y(ext_resp_v_o[4]) );
	BUFX1 U018 ( .A(ext_req_v_i[148]), .Y(local_recv_req) );
	BUFX1 U019 ( .A(local_send_req), .Y(ext_req_v_o[148]) );
	BUFX1 U020 ( .A(ext_resp_v_i[4]), .Y(local_send_resp) );


	MUX21X1 U0(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[24]) ,.Q(int_map_req_v[0]));
	MUX21X1 U1(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[24]) ,.Q(int_map_req_v[1]));
	MUX21X1 U2(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[24]) ,.Q(int_map_req_v[2]));
	MUX21X1 U3(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[24]) ,.Q(int_map_req_v[3]));
	MUX21X1 U4(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[24]) ,.Q(int_map_req_v[4]));
	MUX21X1 U5(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[24]) ,.Q(int_map_req_v[5]));
	MUX21X1 U6(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[24]) ,.Q(int_map_req_v[6]));
	MUX21X1 U7(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[24]) ,.Q(int_map_req_v[7]));
	MUX21X1 U8(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[24]) ,.Q(int_map_req_v[8]));
	MUX21X1 U9(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[24]) ,.Q(int_map_req_v[9]));
	MUX21X1 U10(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[24]) ,.Q(int_map_req_v[10]));
	MUX21X1 U11(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[24]) ,.Q(int_map_req_v[11]));
	MUX21X1 U12(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[24]) ,.Q(int_map_req_v[12]));
	MUX21X1 U13(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[24]) ,.Q(int_map_req_v[13]));
	MUX21X1 U14(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[24]) ,.Q(int_map_req_v[14]));
	MUX21X1 U15(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[24]) ,.Q(int_map_req_v[15]));
	MUX21X1 U16(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[24]) ,.Q(int_map_req_v[16]));
	MUX21X1 U17(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[24]) ,.Q(int_map_req_v[17]));
	MUX21X1 U18(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[24]) ,.Q(int_map_req_v[18]));
	MUX21X1 U19(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[24]) ,.Q(int_map_req_v[19]));
	MUX21X1 U20(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[24]) ,.Q(int_map_req_v[20]));
	MUX21X1 U21(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[24]) ,.Q(int_map_req_v[21]));
	MUX21X1 U22(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[24]) ,.Q(int_map_req_v[22]));
	MUX21X1 U23(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[24]) ,.Q(int_map_req_v[23]));
	MUX21X1 U24(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[24]) ,.Q(int_map_req_v[24]));
	MUX21X1 U25(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[24]) ,.Q(int_map_req_v[25]));
	MUX21X1 U26(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[24]) ,.Q(int_map_req_v[26]));
	MUX21X1 U27(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[24]) ,.Q(int_map_req_v[27]));
	MUX21X1 U28(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[24]) ,.Q(int_map_req_v[28]));
	MUX21X1 U29(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[24]) ,.Q(int_map_req_v[29]));
	MUX21X1 U30(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[24]) ,.Q(int_map_req_v[30]));
	MUX21X1 U31(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[24]) ,.Q(int_map_req_v[31]));
	MUX21X1 U32(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[24]) ,.Q(int_map_req_v[32]));
	MUX21X1 U33(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[24]) ,.Q(int_map_req_v[33]));
	MUX21X1 U34(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[24]) ,.Q(int_map_req_v[34]));
	MUX21X1 U35(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[24]) ,.Q(int_map_req_v[35]));
	MUX21X1 U36(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[24]) ,.Q(int_map_req_v[36]));
	MUX21X1 U37(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[19]) ,.Q(int_map_req_v[37]));
	MUX21X1 U38(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[19]) ,.Q(int_map_req_v[38]));
	MUX21X1 U39(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[19]) ,.Q(int_map_req_v[39]));
	MUX21X1 U40(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[19]) ,.Q(int_map_req_v[40]));
	MUX21X1 U41(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[19]) ,.Q(int_map_req_v[41]));
	MUX21X1 U42(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[19]) ,.Q(int_map_req_v[42]));
	MUX21X1 U43(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[19]) ,.Q(int_map_req_v[43]));
	MUX21X1 U44(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[19]) ,.Q(int_map_req_v[44]));
	MUX21X1 U45(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[19]) ,.Q(int_map_req_v[45]));
	MUX21X1 U46(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[19]) ,.Q(int_map_req_v[46]));
	MUX21X1 U47(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[19]) ,.Q(int_map_req_v[47]));
	MUX21X1 U48(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[19]) ,.Q(int_map_req_v[48]));
	MUX21X1 U49(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[19]) ,.Q(int_map_req_v[49]));
	MUX21X1 U50(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[19]) ,.Q(int_map_req_v[50]));
	MUX21X1 U51(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[19]) ,.Q(int_map_req_v[51]));
	MUX21X1 U52(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[19]) ,.Q(int_map_req_v[52]));
	MUX21X1 U53(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[19]) ,.Q(int_map_req_v[53]));
	MUX21X1 U54(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[19]) ,.Q(int_map_req_v[54]));
	MUX21X1 U55(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[19]) ,.Q(int_map_req_v[55]));
	MUX21X1 U56(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[19]) ,.Q(int_map_req_v[56]));
	MUX21X1 U57(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[19]) ,.Q(int_map_req_v[57]));
	MUX21X1 U58(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[19]) ,.Q(int_map_req_v[58]));
	MUX21X1 U59(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[19]) ,.Q(int_map_req_v[59]));
	MUX21X1 U60(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[19]) ,.Q(int_map_req_v[60]));
	MUX21X1 U61(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[19]) ,.Q(int_map_req_v[61]));
	MUX21X1 U62(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[19]) ,.Q(int_map_req_v[62]));
	MUX21X1 U63(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[19]) ,.Q(int_map_req_v[63]));
	MUX21X1 U64(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[19]) ,.Q(int_map_req_v[64]));
	MUX21X1 U65(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[19]) ,.Q(int_map_req_v[65]));
	MUX21X1 U66(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[19]) ,.Q(int_map_req_v[66]));
	MUX21X1 U67(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[19]) ,.Q(int_map_req_v[67]));
	MUX21X1 U68(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[19]) ,.Q(int_map_req_v[68]));
	MUX21X1 U69(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[19]) ,.Q(int_map_req_v[69]));
	MUX21X1 U70(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[19]) ,.Q(int_map_req_v[70]));
	MUX21X1 U71(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[19]) ,.Q(int_map_req_v[71]));
	MUX21X1 U72(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[19]) ,.Q(int_map_req_v[72]));
	MUX21X1 U73(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[19]) ,.Q(int_map_req_v[73]));
	MUX21X1 U74(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[14]) ,.Q(int_map_req_v[74]));
	MUX21X1 U75(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[14]) ,.Q(int_map_req_v[75]));
	MUX21X1 U76(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[14]) ,.Q(int_map_req_v[76]));
	MUX21X1 U77(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[14]) ,.Q(int_map_req_v[77]));
	MUX21X1 U78(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[14]) ,.Q(int_map_req_v[78]));
	MUX21X1 U79(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[14]) ,.Q(int_map_req_v[79]));
	MUX21X1 U80(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[14]) ,.Q(int_map_req_v[80]));
	MUX21X1 U81(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[14]) ,.Q(int_map_req_v[81]));
	MUX21X1 U82(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[14]) ,.Q(int_map_req_v[82]));
	MUX21X1 U83(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[14]) ,.Q(int_map_req_v[83]));
	MUX21X1 U84(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[14]) ,.Q(int_map_req_v[84]));
	MUX21X1 U85(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[14]) ,.Q(int_map_req_v[85]));
	MUX21X1 U86(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[14]) ,.Q(int_map_req_v[86]));
	MUX21X1 U87(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[14]) ,.Q(int_map_req_v[87]));
	MUX21X1 U88(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[14]) ,.Q(int_map_req_v[88]));
	MUX21X1 U89(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[14]) ,.Q(int_map_req_v[89]));
	MUX21X1 U90(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[14]) ,.Q(int_map_req_v[90]));
	MUX21X1 U91(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[14]) ,.Q(int_map_req_v[91]));
	MUX21X1 U92(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[14]) ,.Q(int_map_req_v[92]));
	MUX21X1 U93(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[14]) ,.Q(int_map_req_v[93]));
	MUX21X1 U94(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[14]) ,.Q(int_map_req_v[94]));
	MUX21X1 U95(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[14]) ,.Q(int_map_req_v[95]));
	MUX21X1 U96(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[14]) ,.Q(int_map_req_v[96]));
	MUX21X1 U97(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[14]) ,.Q(int_map_req_v[97]));
	MUX21X1 U98(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[14]) ,.Q(int_map_req_v[98]));
	MUX21X1 U99(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[14]) ,.Q(int_map_req_v[99]));
	MUX21X1 U100(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[14]) ,.Q(int_map_req_v[100]));
	MUX21X1 U101(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[14]) ,.Q(int_map_req_v[101]));
	MUX21X1 U102(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[14]) ,.Q(int_map_req_v[102]));
	MUX21X1 U103(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[14]) ,.Q(int_map_req_v[103]));
	MUX21X1 U104(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[14]) ,.Q(int_map_req_v[104]));
	MUX21X1 U105(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[14]) ,.Q(int_map_req_v[105]));
	MUX21X1 U106(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[14]) ,.Q(int_map_req_v[106]));
	MUX21X1 U107(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[14]) ,.Q(int_map_req_v[107]));
	MUX21X1 U108(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[14]) ,.Q(int_map_req_v[108]));
	MUX21X1 U109(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[14]) ,.Q(int_map_req_v[109]));
	MUX21X1 U110(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[14]) ,.Q(int_map_req_v[110]));
	MUX21X1 U111(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[9]) ,.Q(int_map_req_v[111]));
	MUX21X1 U112(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[9]) ,.Q(int_map_req_v[112]));
	MUX21X1 U113(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[9]) ,.Q(int_map_req_v[113]));
	MUX21X1 U114(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[9]) ,.Q(int_map_req_v[114]));
	MUX21X1 U115(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[9]) ,.Q(int_map_req_v[115]));
	MUX21X1 U116(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[9]) ,.Q(int_map_req_v[116]));
	MUX21X1 U117(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[9]) ,.Q(int_map_req_v[117]));
	MUX21X1 U118(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[9]) ,.Q(int_map_req_v[118]));
	MUX21X1 U119(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[9]) ,.Q(int_map_req_v[119]));
	MUX21X1 U120(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[9]) ,.Q(int_map_req_v[120]));
	MUX21X1 U121(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[9]) ,.Q(int_map_req_v[121]));
	MUX21X1 U122(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[9]) ,.Q(int_map_req_v[122]));
	MUX21X1 U123(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[9]) ,.Q(int_map_req_v[123]));
	MUX21X1 U124(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[9]) ,.Q(int_map_req_v[124]));
	MUX21X1 U125(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[9]) ,.Q(int_map_req_v[125]));
	MUX21X1 U126(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[9]) ,.Q(int_map_req_v[126]));
	MUX21X1 U127(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[9]) ,.Q(int_map_req_v[127]));
	MUX21X1 U128(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[9]) ,.Q(int_map_req_v[128]));
	MUX21X1 U129(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[9]) ,.Q(int_map_req_v[129]));
	MUX21X1 U130(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[9]) ,.Q(int_map_req_v[130]));
	MUX21X1 U131(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[9]) ,.Q(int_map_req_v[131]));
	MUX21X1 U132(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[9]) ,.Q(int_map_req_v[132]));
	MUX21X1 U133(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[9]) ,.Q(int_map_req_v[133]));
	MUX21X1 U134(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[9]) ,.Q(int_map_req_v[134]));
	MUX21X1 U135(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[9]) ,.Q(int_map_req_v[135]));
	MUX21X1 U136(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[9]) ,.Q(int_map_req_v[136]));
	MUX21X1 U137(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[9]) ,.Q(int_map_req_v[137]));
	MUX21X1 U138(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[9]) ,.Q(int_map_req_v[138]));
	MUX21X1 U139(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[9]) ,.Q(int_map_req_v[139]));
	MUX21X1 U140(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[9]) ,.Q(int_map_req_v[140]));
	MUX21X1 U141(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[9]) ,.Q(int_map_req_v[141]));
	MUX21X1 U142(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[9]) ,.Q(int_map_req_v[142]));
	MUX21X1 U143(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[9]) ,.Q(int_map_req_v[143]));
	MUX21X1 U144(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[9]) ,.Q(int_map_req_v[144]));
	MUX21X1 U145(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[9]) ,.Q(int_map_req_v[145]));
	MUX21X1 U146(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[9]) ,.Q(int_map_req_v[146]));
	MUX21X1 U147(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[9]) ,.Q(int_map_req_v[147]));
	MUX21X1 U01(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[3]), .S(int_route_v[9]) ,.Q(int_resp_v[1]));
	MUX21X1 U02(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[4]), .S(int_route_v[9]) ,.Q(int_resp_v[2]));
	MUX21X1 U03(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[2]), .S(int_route_v[14]) ,.Q(int_resp_v[2]));
	MUX21X1 U04(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[3]), .S(int_route_v[14]) ,.Q(int_resp_v[3]));
	MUX21X1 U05(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[1]), .S(int_route_v[19]) ,.Q(int_resp_v[3]));
	MUX21X1 U06(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[2]), .S(int_route_v[19]) ,.Q(int_resp_v[4]));
	MUX21X1 U07(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[0]), .S(int_route_v[24]) ,.Q(int_resp_v[4]));
	MUX21X1 U08(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[1]), .S(int_route_v[24]) ,.Q(int_resp_v[5]));


	MUX21X1 U148(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[3]) ,.Q(int_map_req_v[148]));
	MUX21X1 U149(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[3]) ,.Q(int_map_req_v[149]));
	MUX21X1 U150(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[3]) ,.Q(int_map_req_v[150]));
	MUX21X1 U151(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[3]) ,.Q(int_map_req_v[151]));
	MUX21X1 U152(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[3]) ,.Q(int_map_req_v[152]));
	MUX21X1 U153(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[3]) ,.Q(int_map_req_v[153]));
	MUX21X1 U154(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[3]) ,.Q(int_map_req_v[154]));
	MUX21X1 U155(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[3]) ,.Q(int_map_req_v[155]));
	MUX21X1 U156(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[3]) ,.Q(int_map_req_v[156]));
	MUX21X1 U157(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[3]) ,.Q(int_map_req_v[157]));
	MUX21X1 U158(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[3]) ,.Q(int_map_req_v[158]));
	MUX21X1 U159(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[3]) ,.Q(int_map_req_v[159]));
	MUX21X1 U160(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[3]) ,.Q(int_map_req_v[160]));
	MUX21X1 U161(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[3]) ,.Q(int_map_req_v[161]));
	MUX21X1 U162(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[3]) ,.Q(int_map_req_v[162]));
	MUX21X1 U163(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[3]) ,.Q(int_map_req_v[163]));
	MUX21X1 U164(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[3]) ,.Q(int_map_req_v[164]));
	MUX21X1 U165(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[3]) ,.Q(int_map_req_v[165]));
	MUX21X1 U166(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[3]) ,.Q(int_map_req_v[166]));
	MUX21X1 U167(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[3]) ,.Q(int_map_req_v[167]));
	MUX21X1 U168(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[3]) ,.Q(int_map_req_v[168]));
	MUX21X1 U169(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[3]) ,.Q(int_map_req_v[169]));
	MUX21X1 U170(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[3]) ,.Q(int_map_req_v[170]));
	MUX21X1 U171(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[3]) ,.Q(int_map_req_v[171]));
	MUX21X1 U172(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[3]) ,.Q(int_map_req_v[172]));
	MUX21X1 U173(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[3]) ,.Q(int_map_req_v[173]));
	MUX21X1 U174(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[3]) ,.Q(int_map_req_v[174]));
	MUX21X1 U175(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[3]) ,.Q(int_map_req_v[175]));
	MUX21X1 U176(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[3]) ,.Q(int_map_req_v[176]));
	MUX21X1 U177(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[3]) ,.Q(int_map_req_v[177]));
	MUX21X1 U178(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[3]) ,.Q(int_map_req_v[178]));
	MUX21X1 U179(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[3]) ,.Q(int_map_req_v[179]));
	MUX21X1 U180(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[3]) ,.Q(int_map_req_v[180]));
	MUX21X1 U181(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[3]) ,.Q(int_map_req_v[181]));
	MUX21X1 U182(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[3]) ,.Q(int_map_req_v[182]));
	MUX21X1 U183(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[3]) ,.Q(int_map_req_v[183]));
	MUX21X1 U184(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[3]) ,.Q(int_map_req_v[184]));
	MUX21X1 U185(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[23]) ,.Q(int_map_req_v[185]));
	MUX21X1 U186(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[23]) ,.Q(int_map_req_v[186]));
	MUX21X1 U187(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[23]) ,.Q(int_map_req_v[187]));
	MUX21X1 U188(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[23]) ,.Q(int_map_req_v[188]));
	MUX21X1 U189(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[23]) ,.Q(int_map_req_v[189]));
	MUX21X1 U190(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[23]) ,.Q(int_map_req_v[190]));
	MUX21X1 U191(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[23]) ,.Q(int_map_req_v[191]));
	MUX21X1 U192(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[23]) ,.Q(int_map_req_v[192]));
	MUX21X1 U193(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[23]) ,.Q(int_map_req_v[193]));
	MUX21X1 U194(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[23]) ,.Q(int_map_req_v[194]));
	MUX21X1 U195(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[23]) ,.Q(int_map_req_v[195]));
	MUX21X1 U196(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[23]) ,.Q(int_map_req_v[196]));
	MUX21X1 U197(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[23]) ,.Q(int_map_req_v[197]));
	MUX21X1 U198(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[23]) ,.Q(int_map_req_v[198]));
	MUX21X1 U199(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[23]) ,.Q(int_map_req_v[199]));
	MUX21X1 U200(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[23]) ,.Q(int_map_req_v[200]));
	MUX21X1 U201(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[23]) ,.Q(int_map_req_v[201]));
	MUX21X1 U202(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[23]) ,.Q(int_map_req_v[202]));
	MUX21X1 U203(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[23]) ,.Q(int_map_req_v[203]));
	MUX21X1 U204(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[23]) ,.Q(int_map_req_v[204]));
	MUX21X1 U205(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[23]) ,.Q(int_map_req_v[205]));
	MUX21X1 U206(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[23]) ,.Q(int_map_req_v[206]));
	MUX21X1 U207(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[23]) ,.Q(int_map_req_v[207]));
	MUX21X1 U208(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[23]) ,.Q(int_map_req_v[208]));
	MUX21X1 U209(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[23]) ,.Q(int_map_req_v[209]));
	MUX21X1 U210(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[23]) ,.Q(int_map_req_v[210]));
	MUX21X1 U211(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[23]) ,.Q(int_map_req_v[211]));
	MUX21X1 U212(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[23]) ,.Q(int_map_req_v[212]));
	MUX21X1 U213(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[23]) ,.Q(int_map_req_v[213]));
	MUX21X1 U214(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[23]) ,.Q(int_map_req_v[214]));
	MUX21X1 U215(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[23]) ,.Q(int_map_req_v[215]));
	MUX21X1 U216(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[23]) ,.Q(int_map_req_v[216]));
	MUX21X1 U217(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[23]) ,.Q(int_map_req_v[217]));
	MUX21X1 U218(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[23]) ,.Q(int_map_req_v[218]));
	MUX21X1 U219(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[23]) ,.Q(int_map_req_v[219]));
	MUX21X1 U220(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[23]) ,.Q(int_map_req_v[220]));
	MUX21X1 U221(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[23]) ,.Q(int_map_req_v[221]));
	MUX21X1 U222(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[18]) ,.Q(int_map_req_v[222]));
	MUX21X1 U223(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[18]) ,.Q(int_map_req_v[223]));
	MUX21X1 U224(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[18]) ,.Q(int_map_req_v[224]));
	MUX21X1 U225(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[18]) ,.Q(int_map_req_v[225]));
	MUX21X1 U226(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[18]) ,.Q(int_map_req_v[226]));
	MUX21X1 U227(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[18]) ,.Q(int_map_req_v[227]));
	MUX21X1 U228(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[18]) ,.Q(int_map_req_v[228]));
	MUX21X1 U229(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[18]) ,.Q(int_map_req_v[229]));
	MUX21X1 U230(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[18]) ,.Q(int_map_req_v[230]));
	MUX21X1 U231(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[18]) ,.Q(int_map_req_v[231]));
	MUX21X1 U232(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[18]) ,.Q(int_map_req_v[232]));
	MUX21X1 U233(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[18]) ,.Q(int_map_req_v[233]));
	MUX21X1 U234(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[18]) ,.Q(int_map_req_v[234]));
	MUX21X1 U235(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[18]) ,.Q(int_map_req_v[235]));
	MUX21X1 U236(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[18]) ,.Q(int_map_req_v[236]));
	MUX21X1 U237(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[18]) ,.Q(int_map_req_v[237]));
	MUX21X1 U238(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[18]) ,.Q(int_map_req_v[238]));
	MUX21X1 U239(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[18]) ,.Q(int_map_req_v[239]));
	MUX21X1 U240(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[18]) ,.Q(int_map_req_v[240]));
	MUX21X1 U241(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[18]) ,.Q(int_map_req_v[241]));
	MUX21X1 U242(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[18]) ,.Q(int_map_req_v[242]));
	MUX21X1 U243(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[18]) ,.Q(int_map_req_v[243]));
	MUX21X1 U244(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[18]) ,.Q(int_map_req_v[244]));
	MUX21X1 U245(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[18]) ,.Q(int_map_req_v[245]));
	MUX21X1 U246(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[18]) ,.Q(int_map_req_v[246]));
	MUX21X1 U247(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[18]) ,.Q(int_map_req_v[247]));
	MUX21X1 U248(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[18]) ,.Q(int_map_req_v[248]));
	MUX21X1 U249(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[18]) ,.Q(int_map_req_v[249]));
	MUX21X1 U250(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[18]) ,.Q(int_map_req_v[250]));
	MUX21X1 U251(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[18]) ,.Q(int_map_req_v[251]));
	MUX21X1 U252(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[18]) ,.Q(int_map_req_v[252]));
	MUX21X1 U253(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[18]) ,.Q(int_map_req_v[253]));
	MUX21X1 U254(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[18]) ,.Q(int_map_req_v[254]));
	MUX21X1 U255(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[18]) ,.Q(int_map_req_v[255]));
	MUX21X1 U256(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[18]) ,.Q(int_map_req_v[256]));
	MUX21X1 U257(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[18]) ,.Q(int_map_req_v[257]));
	MUX21X1 U258(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[18]) ,.Q(int_map_req_v[258]));
	MUX21X1 U259(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[13]) ,.Q(int_map_req_v[259]));
	MUX21X1 U260(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[13]) ,.Q(int_map_req_v[260]));
	MUX21X1 U261(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[13]) ,.Q(int_map_req_v[261]));
	MUX21X1 U262(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[13]) ,.Q(int_map_req_v[262]));
	MUX21X1 U263(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[13]) ,.Q(int_map_req_v[263]));
	MUX21X1 U264(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[13]) ,.Q(int_map_req_v[264]));
	MUX21X1 U265(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[13]) ,.Q(int_map_req_v[265]));
	MUX21X1 U266(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[13]) ,.Q(int_map_req_v[266]));
	MUX21X1 U267(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[13]) ,.Q(int_map_req_v[267]));
	MUX21X1 U268(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[13]) ,.Q(int_map_req_v[268]));
	MUX21X1 U269(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[13]) ,.Q(int_map_req_v[269]));
	MUX21X1 U270(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[13]) ,.Q(int_map_req_v[270]));
	MUX21X1 U271(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[13]) ,.Q(int_map_req_v[271]));
	MUX21X1 U272(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[13]) ,.Q(int_map_req_v[272]));
	MUX21X1 U273(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[13]) ,.Q(int_map_req_v[273]));
	MUX21X1 U274(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[13]) ,.Q(int_map_req_v[274]));
	MUX21X1 U275(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[13]) ,.Q(int_map_req_v[275]));
	MUX21X1 U276(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[13]) ,.Q(int_map_req_v[276]));
	MUX21X1 U277(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[13]) ,.Q(int_map_req_v[277]));
	MUX21X1 U278(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[13]) ,.Q(int_map_req_v[278]));
	MUX21X1 U279(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[13]) ,.Q(int_map_req_v[279]));
	MUX21X1 U280(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[13]) ,.Q(int_map_req_v[280]));
	MUX21X1 U281(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[13]) ,.Q(int_map_req_v[281]));
	MUX21X1 U282(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[13]) ,.Q(int_map_req_v[282]));
	MUX21X1 U283(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[13]) ,.Q(int_map_req_v[283]));
	MUX21X1 U284(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[13]) ,.Q(int_map_req_v[284]));
	MUX21X1 U285(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[13]) ,.Q(int_map_req_v[285]));
	MUX21X1 U286(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[13]) ,.Q(int_map_req_v[286]));
	MUX21X1 U287(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[13]) ,.Q(int_map_req_v[287]));
	MUX21X1 U288(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[13]) ,.Q(int_map_req_v[288]));
	MUX21X1 U289(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[13]) ,.Q(int_map_req_v[289]));
	MUX21X1 U290(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[13]) ,.Q(int_map_req_v[290]));
	MUX21X1 U291(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[13]) ,.Q(int_map_req_v[291]));
	MUX21X1 U292(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[13]) ,.Q(int_map_req_v[292]));
	MUX21X1 U293(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[13]) ,.Q(int_map_req_v[293]));
	MUX21X1 U294(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[13]) ,.Q(int_map_req_v[294]));
	MUX21X1 U295(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[13]) ,.Q(int_map_req_v[295]));
	MUX21X1 U09(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[7]), .S(int_route_v[13]) ,.Q(int_resp_v[2]));
	MUX21X1 U10(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[8]), .S(int_route_v[13]) ,.Q(int_resp_v[3]));
	MUX21X1 U11(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[6]), .S(int_route_v[18]) ,.Q(int_resp_v[3]));
	MUX21X1 U12(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[7]), .S(int_route_v[18]) ,.Q(int_resp_v[4]));
	MUX21X1 U13(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[4]));
	MUX21X1 U14(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[2]), .S(int_route_v[6]) ,.Q(int_resp_v[5]));
	MUX21X1 U15(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[0]), .S(int_route_v[4]) ,.Q(int_resp_v[0]));
	MUX21X1 U16(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));


	MUX21X1 U296(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[7]) ,.Q(int_map_req_v[296]));
	MUX21X1 U297(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[7]) ,.Q(int_map_req_v[297]));
	MUX21X1 U298(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[7]) ,.Q(int_map_req_v[298]));
	MUX21X1 U299(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[7]) ,.Q(int_map_req_v[299]));
	MUX21X1 U300(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[7]) ,.Q(int_map_req_v[300]));
	MUX21X1 U301(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[7]) ,.Q(int_map_req_v[301]));
	MUX21X1 U302(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[7]) ,.Q(int_map_req_v[302]));
	MUX21X1 U303(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[7]) ,.Q(int_map_req_v[303]));
	MUX21X1 U304(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[7]) ,.Q(int_map_req_v[304]));
	MUX21X1 U305(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[7]) ,.Q(int_map_req_v[305]));
	MUX21X1 U306(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[7]) ,.Q(int_map_req_v[306]));
	MUX21X1 U307(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[7]) ,.Q(int_map_req_v[307]));
	MUX21X1 U308(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[7]) ,.Q(int_map_req_v[308]));
	MUX21X1 U309(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[7]) ,.Q(int_map_req_v[309]));
	MUX21X1 U310(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[7]) ,.Q(int_map_req_v[310]));
	MUX21X1 U311(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[7]) ,.Q(int_map_req_v[311]));
	MUX21X1 U312(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[7]) ,.Q(int_map_req_v[312]));
	MUX21X1 U313(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[7]) ,.Q(int_map_req_v[313]));
	MUX21X1 U314(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[7]) ,.Q(int_map_req_v[314]));
	MUX21X1 U315(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[7]) ,.Q(int_map_req_v[315]));
	MUX21X1 U316(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[7]) ,.Q(int_map_req_v[316]));
	MUX21X1 U317(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[7]) ,.Q(int_map_req_v[317]));
	MUX21X1 U318(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[7]) ,.Q(int_map_req_v[318]));
	MUX21X1 U319(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[7]) ,.Q(int_map_req_v[319]));
	MUX21X1 U320(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[7]) ,.Q(int_map_req_v[320]));
	MUX21X1 U321(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[7]) ,.Q(int_map_req_v[321]));
	MUX21X1 U322(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[7]) ,.Q(int_map_req_v[322]));
	MUX21X1 U323(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[7]) ,.Q(int_map_req_v[323]));
	MUX21X1 U324(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[7]) ,.Q(int_map_req_v[324]));
	MUX21X1 U325(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[7]) ,.Q(int_map_req_v[325]));
	MUX21X1 U326(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[7]) ,.Q(int_map_req_v[326]));
	MUX21X1 U327(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[7]) ,.Q(int_map_req_v[327]));
	MUX21X1 U328(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[7]) ,.Q(int_map_req_v[328]));
	MUX21X1 U329(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[7]) ,.Q(int_map_req_v[329]));
	MUX21X1 U330(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[7]) ,.Q(int_map_req_v[330]));
	MUX21X1 U331(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[7]) ,.Q(int_map_req_v[331]));
	MUX21X1 U332(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[7]) ,.Q(int_map_req_v[332]));
	MUX21X1 U333(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[2]) ,.Q(int_map_req_v[333]));
	MUX21X1 U334(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[2]) ,.Q(int_map_req_v[334]));
	MUX21X1 U335(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[2]) ,.Q(int_map_req_v[335]));
	MUX21X1 U336(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[2]) ,.Q(int_map_req_v[336]));
	MUX21X1 U337(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[2]) ,.Q(int_map_req_v[337]));
	MUX21X1 U338(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[2]) ,.Q(int_map_req_v[338]));
	MUX21X1 U339(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[2]) ,.Q(int_map_req_v[339]));
	MUX21X1 U340(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[2]) ,.Q(int_map_req_v[340]));
	MUX21X1 U341(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[2]) ,.Q(int_map_req_v[341]));
	MUX21X1 U342(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[2]) ,.Q(int_map_req_v[342]));
	MUX21X1 U343(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[2]) ,.Q(int_map_req_v[343]));
	MUX21X1 U344(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[2]) ,.Q(int_map_req_v[344]));
	MUX21X1 U345(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[2]) ,.Q(int_map_req_v[345]));
	MUX21X1 U346(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[2]) ,.Q(int_map_req_v[346]));
	MUX21X1 U347(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[2]) ,.Q(int_map_req_v[347]));
	MUX21X1 U348(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[2]) ,.Q(int_map_req_v[348]));
	MUX21X1 U349(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[2]) ,.Q(int_map_req_v[349]));
	MUX21X1 U350(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[2]) ,.Q(int_map_req_v[350]));
	MUX21X1 U351(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[2]) ,.Q(int_map_req_v[351]));
	MUX21X1 U352(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[2]) ,.Q(int_map_req_v[352]));
	MUX21X1 U353(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[2]) ,.Q(int_map_req_v[353]));
	MUX21X1 U354(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[2]) ,.Q(int_map_req_v[354]));
	MUX21X1 U355(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[2]) ,.Q(int_map_req_v[355]));
	MUX21X1 U356(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[2]) ,.Q(int_map_req_v[356]));
	MUX21X1 U357(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[2]) ,.Q(int_map_req_v[357]));
	MUX21X1 U358(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[2]) ,.Q(int_map_req_v[358]));
	MUX21X1 U359(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[2]) ,.Q(int_map_req_v[359]));
	MUX21X1 U360(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[2]) ,.Q(int_map_req_v[360]));
	MUX21X1 U361(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[2]) ,.Q(int_map_req_v[361]));
	MUX21X1 U362(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[2]) ,.Q(int_map_req_v[362]));
	MUX21X1 U363(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[2]) ,.Q(int_map_req_v[363]));
	MUX21X1 U364(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[2]) ,.Q(int_map_req_v[364]));
	MUX21X1 U365(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[2]) ,.Q(int_map_req_v[365]));
	MUX21X1 U366(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[2]) ,.Q(int_map_req_v[366]));
	MUX21X1 U367(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[2]) ,.Q(int_map_req_v[367]));
	MUX21X1 U368(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[2]) ,.Q(int_map_req_v[368]));
	MUX21X1 U369(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[2]) ,.Q(int_map_req_v[369]));
	MUX21X1 U370(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[22]) ,.Q(int_map_req_v[370]));
	MUX21X1 U371(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[22]) ,.Q(int_map_req_v[371]));
	MUX21X1 U372(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[22]) ,.Q(int_map_req_v[372]));
	MUX21X1 U373(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[22]) ,.Q(int_map_req_v[373]));
	MUX21X1 U374(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[22]) ,.Q(int_map_req_v[374]));
	MUX21X1 U375(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[22]) ,.Q(int_map_req_v[375]));
	MUX21X1 U376(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[22]) ,.Q(int_map_req_v[376]));
	MUX21X1 U377(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[22]) ,.Q(int_map_req_v[377]));
	MUX21X1 U378(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[22]) ,.Q(int_map_req_v[378]));
	MUX21X1 U379(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[22]) ,.Q(int_map_req_v[379]));
	MUX21X1 U380(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[22]) ,.Q(int_map_req_v[380]));
	MUX21X1 U381(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[22]) ,.Q(int_map_req_v[381]));
	MUX21X1 U382(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[22]) ,.Q(int_map_req_v[382]));
	MUX21X1 U383(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[22]) ,.Q(int_map_req_v[383]));
	MUX21X1 U384(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[22]) ,.Q(int_map_req_v[384]));
	MUX21X1 U385(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[22]) ,.Q(int_map_req_v[385]));
	MUX21X1 U386(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[22]) ,.Q(int_map_req_v[386]));
	MUX21X1 U387(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[22]) ,.Q(int_map_req_v[387]));
	MUX21X1 U388(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[22]) ,.Q(int_map_req_v[388]));
	MUX21X1 U389(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[22]) ,.Q(int_map_req_v[389]));
	MUX21X1 U390(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[22]) ,.Q(int_map_req_v[390]));
	MUX21X1 U391(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[22]) ,.Q(int_map_req_v[391]));
	MUX21X1 U392(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[22]) ,.Q(int_map_req_v[392]));
	MUX21X1 U393(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[22]) ,.Q(int_map_req_v[393]));
	MUX21X1 U394(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[22]) ,.Q(int_map_req_v[394]));
	MUX21X1 U395(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[22]) ,.Q(int_map_req_v[395]));
	MUX21X1 U396(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[22]) ,.Q(int_map_req_v[396]));
	MUX21X1 U397(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[22]) ,.Q(int_map_req_v[397]));
	MUX21X1 U398(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[22]) ,.Q(int_map_req_v[398]));
	MUX21X1 U399(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[22]) ,.Q(int_map_req_v[399]));
	MUX21X1 U400(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[22]) ,.Q(int_map_req_v[400]));
	MUX21X1 U401(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[22]) ,.Q(int_map_req_v[401]));
	MUX21X1 U402(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[22]) ,.Q(int_map_req_v[402]));
	MUX21X1 U403(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[22]) ,.Q(int_map_req_v[403]));
	MUX21X1 U404(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[22]) ,.Q(int_map_req_v[404]));
	MUX21X1 U405(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[22]) ,.Q(int_map_req_v[405]));
	MUX21X1 U406(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[22]) ,.Q(int_map_req_v[406]));
	MUX21X1 U407(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[17]) ,.Q(int_map_req_v[407]));
	MUX21X1 U408(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[17]) ,.Q(int_map_req_v[408]));
	MUX21X1 U409(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[17]) ,.Q(int_map_req_v[409]));
	MUX21X1 U410(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[17]) ,.Q(int_map_req_v[410]));
	MUX21X1 U411(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[17]) ,.Q(int_map_req_v[411]));
	MUX21X1 U412(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[17]) ,.Q(int_map_req_v[412]));
	MUX21X1 U413(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[17]) ,.Q(int_map_req_v[413]));
	MUX21X1 U414(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[17]) ,.Q(int_map_req_v[414]));
	MUX21X1 U415(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[17]) ,.Q(int_map_req_v[415]));
	MUX21X1 U416(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[17]) ,.Q(int_map_req_v[416]));
	MUX21X1 U417(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[17]) ,.Q(int_map_req_v[417]));
	MUX21X1 U418(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[17]) ,.Q(int_map_req_v[418]));
	MUX21X1 U419(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[17]) ,.Q(int_map_req_v[419]));
	MUX21X1 U420(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[17]) ,.Q(int_map_req_v[420]));
	MUX21X1 U421(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[17]) ,.Q(int_map_req_v[421]));
	MUX21X1 U422(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[17]) ,.Q(int_map_req_v[422]));
	MUX21X1 U423(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[17]) ,.Q(int_map_req_v[423]));
	MUX21X1 U424(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[17]) ,.Q(int_map_req_v[424]));
	MUX21X1 U425(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[17]) ,.Q(int_map_req_v[425]));
	MUX21X1 U426(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[17]) ,.Q(int_map_req_v[426]));
	MUX21X1 U427(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[17]) ,.Q(int_map_req_v[427]));
	MUX21X1 U428(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[17]) ,.Q(int_map_req_v[428]));
	MUX21X1 U429(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[17]) ,.Q(int_map_req_v[429]));
	MUX21X1 U430(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[17]) ,.Q(int_map_req_v[430]));
	MUX21X1 U431(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[17]) ,.Q(int_map_req_v[431]));
	MUX21X1 U432(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[17]) ,.Q(int_map_req_v[432]));
	MUX21X1 U433(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[17]) ,.Q(int_map_req_v[433]));
	MUX21X1 U434(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[17]) ,.Q(int_map_req_v[434]));
	MUX21X1 U435(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[17]) ,.Q(int_map_req_v[435]));
	MUX21X1 U436(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[17]) ,.Q(int_map_req_v[436]));
	MUX21X1 U437(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[17]) ,.Q(int_map_req_v[437]));
	MUX21X1 U438(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[17]) ,.Q(int_map_req_v[438]));
	MUX21X1 U439(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[17]) ,.Q(int_map_req_v[439]));
	MUX21X1 U440(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[17]) ,.Q(int_map_req_v[440]));
	MUX21X1 U441(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[17]) ,.Q(int_map_req_v[441]));
	MUX21X1 U442(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[17]) ,.Q(int_map_req_v[442]));
	MUX21X1 U443(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[17]) ,.Q(int_map_req_v[443]));
	MUX21X1 U17(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[11]), .S(int_route_v[17]) ,.Q(int_resp_v[3]));
	MUX21X1 U18(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[12]), .S(int_route_v[17]) ,.Q(int_resp_v[4]));
	MUX21X1 U19(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[10]), .S(int_route_v[22]) ,.Q(int_resp_v[4]));
	MUX21X1 U20(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[11]), .S(int_route_v[22]) ,.Q(int_resp_v[5]));
	MUX21X1 U21(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[9]), .S(int_route_v[2]) ,.Q(int_resp_v[0]));
	MUX21X1 U22(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[10]), .S(int_route_v[2]) ,.Q(int_resp_v[1]));
	MUX21X1 U23(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[8]), .S(int_route_v[7]) ,.Q(int_resp_v[1]));
	MUX21X1 U24(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[9]), .S(int_route_v[7]) ,.Q(int_resp_v[2]));

	MUX21X1 U444(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[11]) ,.Q(int_map_req_v[444]));
	MUX21X1 U445(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[11]) ,.Q(int_map_req_v[445]));
	MUX21X1 U446(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[11]) ,.Q(int_map_req_v[446]));
	MUX21X1 U447(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[11]) ,.Q(int_map_req_v[447]));
	MUX21X1 U448(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[11]) ,.Q(int_map_req_v[448]));
	MUX21X1 U449(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[11]) ,.Q(int_map_req_v[449]));
	MUX21X1 U450(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[11]) ,.Q(int_map_req_v[450]));
	MUX21X1 U451(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[11]) ,.Q(int_map_req_v[451]));
	MUX21X1 U452(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[11]) ,.Q(int_map_req_v[452]));
	MUX21X1 U453(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[11]) ,.Q(int_map_req_v[453]));
	MUX21X1 U454(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[11]) ,.Q(int_map_req_v[454]));
	MUX21X1 U455(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[11]) ,.Q(int_map_req_v[455]));
	MUX21X1 U456(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[11]) ,.Q(int_map_req_v[456]));
	MUX21X1 U457(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[11]) ,.Q(int_map_req_v[457]));
	MUX21X1 U458(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[11]) ,.Q(int_map_req_v[458]));
	MUX21X1 U459(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[11]) ,.Q(int_map_req_v[459]));
	MUX21X1 U460(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[11]) ,.Q(int_map_req_v[460]));
	MUX21X1 U461(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[11]) ,.Q(int_map_req_v[461]));
	MUX21X1 U462(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[11]) ,.Q(int_map_req_v[462]));
	MUX21X1 U463(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[11]) ,.Q(int_map_req_v[463]));
	MUX21X1 U464(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[11]) ,.Q(int_map_req_v[464]));
	MUX21X1 U465(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[11]) ,.Q(int_map_req_v[465]));
	MUX21X1 U466(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[11]) ,.Q(int_map_req_v[466]));
	MUX21X1 U467(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[11]) ,.Q(int_map_req_v[467]));
	MUX21X1 U468(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[11]) ,.Q(int_map_req_v[468]));
	MUX21X1 U469(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[11]) ,.Q(int_map_req_v[469]));
	MUX21X1 U470(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[11]) ,.Q(int_map_req_v[470]));
	MUX21X1 U471(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[11]) ,.Q(int_map_req_v[471]));
	MUX21X1 U472(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[11]) ,.Q(int_map_req_v[472]));
	MUX21X1 U473(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[11]) ,.Q(int_map_req_v[473]));
	MUX21X1 U474(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[11]) ,.Q(int_map_req_v[474]));
	MUX21X1 U475(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[11]) ,.Q(int_map_req_v[475]));
	MUX21X1 U476(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[11]) ,.Q(int_map_req_v[476]));
	MUX21X1 U477(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[11]) ,.Q(int_map_req_v[477]));
	MUX21X1 U478(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[11]) ,.Q(int_map_req_v[478]));
	MUX21X1 U479(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[11]) ,.Q(int_map_req_v[479]));
	MUX21X1 U480(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[11]) ,.Q(int_map_req_v[480]));
	MUX21X1 U481(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[6]) ,.Q(int_map_req_v[481]));
	MUX21X1 U482(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[6]) ,.Q(int_map_req_v[482]));
	MUX21X1 U483(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[6]) ,.Q(int_map_req_v[483]));
	MUX21X1 U484(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[6]) ,.Q(int_map_req_v[484]));
	MUX21X1 U485(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[6]) ,.Q(int_map_req_v[485]));
	MUX21X1 U486(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[6]) ,.Q(int_map_req_v[486]));
	MUX21X1 U487(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[6]) ,.Q(int_map_req_v[487]));
	MUX21X1 U488(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[6]) ,.Q(int_map_req_v[488]));
	MUX21X1 U489(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[6]) ,.Q(int_map_req_v[489]));
	MUX21X1 U490(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[6]) ,.Q(int_map_req_v[490]));
	MUX21X1 U491(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[6]) ,.Q(int_map_req_v[491]));
	MUX21X1 U492(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[6]) ,.Q(int_map_req_v[492]));
	MUX21X1 U493(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[6]) ,.Q(int_map_req_v[493]));
	MUX21X1 U494(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[6]) ,.Q(int_map_req_v[494]));
	MUX21X1 U495(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[6]) ,.Q(int_map_req_v[495]));
	MUX21X1 U496(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[6]) ,.Q(int_map_req_v[496]));
	MUX21X1 U497(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[6]) ,.Q(int_map_req_v[497]));
	MUX21X1 U498(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[6]) ,.Q(int_map_req_v[498]));
	MUX21X1 U499(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[6]) ,.Q(int_map_req_v[499]));
	MUX21X1 U500(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[6]) ,.Q(int_map_req_v[500]));
	MUX21X1 U501(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[6]) ,.Q(int_map_req_v[501]));
	MUX21X1 U502(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[6]) ,.Q(int_map_req_v[502]));
	MUX21X1 U503(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[6]) ,.Q(int_map_req_v[503]));
	MUX21X1 U504(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[6]) ,.Q(int_map_req_v[504]));
	MUX21X1 U505(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[6]) ,.Q(int_map_req_v[505]));
	MUX21X1 U506(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[6]) ,.Q(int_map_req_v[506]));
	MUX21X1 U507(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[6]) ,.Q(int_map_req_v[507]));
	MUX21X1 U508(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[6]) ,.Q(int_map_req_v[508]));
	MUX21X1 U509(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[6]) ,.Q(int_map_req_v[509]));
	MUX21X1 U510(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[6]) ,.Q(int_map_req_v[510]));
	MUX21X1 U511(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[6]) ,.Q(int_map_req_v[511]));
	MUX21X1 U512(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[6]) ,.Q(int_map_req_v[512]));
	MUX21X1 U513(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[6]) ,.Q(int_map_req_v[513]));
	MUX21X1 U514(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[6]) ,.Q(int_map_req_v[514]));
	MUX21X1 U515(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[6]) ,.Q(int_map_req_v[515]));
	MUX21X1 U516(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[6]) ,.Q(int_map_req_v[516]));
	MUX21X1 U517(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[6]) ,.Q(int_map_req_v[517]));
	MUX21X1 U518(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[1]) ,.Q(int_map_req_v[518]));
	MUX21X1 U519(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[1]) ,.Q(int_map_req_v[519]));
	MUX21X1 U520(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[1]) ,.Q(int_map_req_v[520]));
	MUX21X1 U521(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[1]) ,.Q(int_map_req_v[521]));
	MUX21X1 U522(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[1]) ,.Q(int_map_req_v[522]));
	MUX21X1 U523(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[1]) ,.Q(int_map_req_v[523]));
	MUX21X1 U524(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[1]) ,.Q(int_map_req_v[524]));
	MUX21X1 U525(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[1]) ,.Q(int_map_req_v[525]));
	MUX21X1 U526(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[1]) ,.Q(int_map_req_v[526]));
	MUX21X1 U527(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[1]) ,.Q(int_map_req_v[527]));
	MUX21X1 U528(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[1]) ,.Q(int_map_req_v[528]));
	MUX21X1 U529(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[1]) ,.Q(int_map_req_v[529]));
	MUX21X1 U530(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[1]) ,.Q(int_map_req_v[530]));
	MUX21X1 U531(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[1]) ,.Q(int_map_req_v[531]));
	MUX21X1 U532(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[1]) ,.Q(int_map_req_v[532]));
	MUX21X1 U533(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[1]) ,.Q(int_map_req_v[533]));
	MUX21X1 U534(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[1]) ,.Q(int_map_req_v[534]));
	MUX21X1 U535(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[1]) ,.Q(int_map_req_v[535]));
	MUX21X1 U536(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[1]) ,.Q(int_map_req_v[536]));
	MUX21X1 U537(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[1]) ,.Q(int_map_req_v[537]));
	MUX21X1 U538(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[1]) ,.Q(int_map_req_v[538]));
	MUX21X1 U539(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[1]) ,.Q(int_map_req_v[539]));
	MUX21X1 U540(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[1]) ,.Q(int_map_req_v[540]));
	MUX21X1 U541(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[1]) ,.Q(int_map_req_v[541]));
	MUX21X1 U542(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[1]) ,.Q(int_map_req_v[542]));
	MUX21X1 U543(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[1]) ,.Q(int_map_req_v[543]));
	MUX21X1 U544(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[1]) ,.Q(int_map_req_v[544]));
	MUX21X1 U545(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[1]) ,.Q(int_map_req_v[545]));
	MUX21X1 U546(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[1]) ,.Q(int_map_req_v[546]));
	MUX21X1 U547(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[1]) ,.Q(int_map_req_v[547]));
	MUX21X1 U548(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[1]) ,.Q(int_map_req_v[548]));
	MUX21X1 U549(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[1]) ,.Q(int_map_req_v[549]));
	MUX21X1 U550(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[1]) ,.Q(int_map_req_v[550]));
	MUX21X1 U551(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[1]) ,.Q(int_map_req_v[551]));
	MUX21X1 U552(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[1]) ,.Q(int_map_req_v[552]));
	MUX21X1 U553(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[1]) ,.Q(int_map_req_v[553]));
	MUX21X1 U554(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[1]) ,.Q(int_map_req_v[554]));
	MUX21X1 U555(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[21]) ,.Q(int_map_req_v[555]));
	MUX21X1 U556(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[21]) ,.Q(int_map_req_v[556]));
	MUX21X1 U557(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[21]) ,.Q(int_map_req_v[557]));
	MUX21X1 U558(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[21]) ,.Q(int_map_req_v[558]));
	MUX21X1 U559(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[21]) ,.Q(int_map_req_v[559]));
	MUX21X1 U560(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[21]) ,.Q(int_map_req_v[560]));
	MUX21X1 U561(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[21]) ,.Q(int_map_req_v[561]));
	MUX21X1 U562(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[21]) ,.Q(int_map_req_v[562]));
	MUX21X1 U563(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[21]) ,.Q(int_map_req_v[563]));
	MUX21X1 U564(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[21]) ,.Q(int_map_req_v[564]));
	MUX21X1 U565(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[21]) ,.Q(int_map_req_v[565]));
	MUX21X1 U566(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[21]) ,.Q(int_map_req_v[566]));
	MUX21X1 U567(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[21]) ,.Q(int_map_req_v[567]));
	MUX21X1 U568(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[21]) ,.Q(int_map_req_v[568]));
	MUX21X1 U569(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[21]) ,.Q(int_map_req_v[569]));
	MUX21X1 U570(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[21]) ,.Q(int_map_req_v[570]));
	MUX21X1 U571(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[21]) ,.Q(int_map_req_v[571]));
	MUX21X1 U572(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[21]) ,.Q(int_map_req_v[572]));
	MUX21X1 U573(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[21]) ,.Q(int_map_req_v[573]));
	MUX21X1 U574(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[21]) ,.Q(int_map_req_v[574]));
	MUX21X1 U575(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[21]) ,.Q(int_map_req_v[575]));
	MUX21X1 U576(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[21]) ,.Q(int_map_req_v[576]));
	MUX21X1 U577(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[21]) ,.Q(int_map_req_v[577]));
	MUX21X1 U578(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[21]) ,.Q(int_map_req_v[578]));
	MUX21X1 U579(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[21]) ,.Q(int_map_req_v[579]));
	MUX21X1 U580(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[21]) ,.Q(int_map_req_v[580]));
	MUX21X1 U581(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[21]) ,.Q(int_map_req_v[581]));
	MUX21X1 U582(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[21]) ,.Q(int_map_req_v[582]));
	MUX21X1 U583(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[21]) ,.Q(int_map_req_v[583]));
	MUX21X1 U584(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[21]) ,.Q(int_map_req_v[584]));
	MUX21X1 U585(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[21]) ,.Q(int_map_req_v[585]));
	MUX21X1 U586(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[21]) ,.Q(int_map_req_v[586]));
	MUX21X1 U587(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[21]) ,.Q(int_map_req_v[587]));
	MUX21X1 U588(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[21]) ,.Q(int_map_req_v[588]));
	MUX21X1 U589(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[21]) ,.Q(int_map_req_v[589]));
	MUX21X1 U590(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[21]) ,.Q(int_map_req_v[590]));
	MUX21X1 U591(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[21]) ,.Q(int_map_req_v[591]));
	MUX21X1 U25(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[15]), .S(int_route_v[21]) ,.Q(int_resp_v[4]));
	MUX21X1 U26(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[16]), .S(int_route_v[21]) ,.Q(int_resp_v[5]));
	MUX21X1 U27(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[14]), .S(int_route_v[1]) ,.Q(int_resp_v[0]));
	MUX21X1 U28(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[15]), .S(int_route_v[1]) ,.Q(int_resp_v[1]));
	MUX21X1 U29(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[13]), .S(int_route_v[6]) ,.Q(int_resp_v[1]));
	MUX21X1 U30(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[14]), .S(int_route_v[6]) ,.Q(int_resp_v[2]));
	MUX21X1 U31(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[12]), .S(int_route_v[11]) ,.Q(int_resp_v[2]));
	MUX21X1 U32(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[13]), .S(int_route_v[11]) ,.Q(int_resp_v[3]));



	MUX21X1 U592(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[15]) ,.Q(int_map_req_v[592]));
	MUX21X1 U593(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[15]) ,.Q(int_map_req_v[593]));
	MUX21X1 U594(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[15]) ,.Q(int_map_req_v[594]));
	MUX21X1 U595(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[15]) ,.Q(int_map_req_v[595]));
	MUX21X1 U596(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[15]) ,.Q(int_map_req_v[596]));
	MUX21X1 U597(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[15]) ,.Q(int_map_req_v[597]));
	MUX21X1 U598(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[15]) ,.Q(int_map_req_v[598]));
	MUX21X1 U599(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[15]) ,.Q(int_map_req_v[599]));
	MUX21X1 U600(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[15]) ,.Q(int_map_req_v[600]));
	MUX21X1 U601(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[15]) ,.Q(int_map_req_v[601]));
	MUX21X1 U602(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[15]) ,.Q(int_map_req_v[602]));
	MUX21X1 U603(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[15]) ,.Q(int_map_req_v[603]));
	MUX21X1 U604(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[15]) ,.Q(int_map_req_v[604]));
	MUX21X1 U605(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[15]) ,.Q(int_map_req_v[605]));
	MUX21X1 U606(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[15]) ,.Q(int_map_req_v[606]));
	MUX21X1 U607(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[15]) ,.Q(int_map_req_v[607]));
	MUX21X1 U608(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[15]) ,.Q(int_map_req_v[608]));
	MUX21X1 U609(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[15]) ,.Q(int_map_req_v[609]));
	MUX21X1 U610(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[15]) ,.Q(int_map_req_v[610]));
	MUX21X1 U611(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[15]) ,.Q(int_map_req_v[611]));
	MUX21X1 U612(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[15]) ,.Q(int_map_req_v[612]));
	MUX21X1 U613(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[15]) ,.Q(int_map_req_v[613]));
	MUX21X1 U614(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[15]) ,.Q(int_map_req_v[614]));
	MUX21X1 U615(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[15]) ,.Q(int_map_req_v[615]));
	MUX21X1 U616(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[15]) ,.Q(int_map_req_v[616]));
	MUX21X1 U617(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[15]) ,.Q(int_map_req_v[617]));
	MUX21X1 U618(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[15]) ,.Q(int_map_req_v[618]));
	MUX21X1 U619(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[15]) ,.Q(int_map_req_v[619]));
	MUX21X1 U620(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[15]) ,.Q(int_map_req_v[620]));
	MUX21X1 U621(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[15]) ,.Q(int_map_req_v[621]));
	MUX21X1 U622(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[15]) ,.Q(int_map_req_v[622]));
	MUX21X1 U623(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[15]) ,.Q(int_map_req_v[623]));
	MUX21X1 U624(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[15]) ,.Q(int_map_req_v[624]));
	MUX21X1 U625(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[15]) ,.Q(int_map_req_v[625]));
	MUX21X1 U626(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[15]) ,.Q(int_map_req_v[626]));
	MUX21X1 U627(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[15]) ,.Q(int_map_req_v[627]));
	MUX21X1 U628(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[15]) ,.Q(int_map_req_v[628]));
	MUX21X1 U629(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[10]) ,.Q(int_map_req_v[629]));
	MUX21X1 U630(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[10]) ,.Q(int_map_req_v[630]));
	MUX21X1 U631(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[10]) ,.Q(int_map_req_v[631]));
	MUX21X1 U632(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[10]) ,.Q(int_map_req_v[632]));
	MUX21X1 U633(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[10]) ,.Q(int_map_req_v[633]));
	MUX21X1 U634(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[10]) ,.Q(int_map_req_v[634]));
	MUX21X1 U635(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[10]) ,.Q(int_map_req_v[635]));
	MUX21X1 U636(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[10]) ,.Q(int_map_req_v[636]));
	MUX21X1 U637(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[10]) ,.Q(int_map_req_v[637]));
	MUX21X1 U638(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[10]) ,.Q(int_map_req_v[638]));
	MUX21X1 U639(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[10]) ,.Q(int_map_req_v[639]));
	MUX21X1 U640(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[10]) ,.Q(int_map_req_v[640]));
	MUX21X1 U641(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[10]) ,.Q(int_map_req_v[641]));
	MUX21X1 U642(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[10]) ,.Q(int_map_req_v[642]));
	MUX21X1 U643(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[10]) ,.Q(int_map_req_v[643]));
	MUX21X1 U644(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[10]) ,.Q(int_map_req_v[644]));
	MUX21X1 U645(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[10]) ,.Q(int_map_req_v[645]));
	MUX21X1 U646(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[10]) ,.Q(int_map_req_v[646]));
	MUX21X1 U647(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[10]) ,.Q(int_map_req_v[647]));
	MUX21X1 U648(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[10]) ,.Q(int_map_req_v[648]));
	MUX21X1 U649(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[10]) ,.Q(int_map_req_v[649]));
	MUX21X1 U650(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[10]) ,.Q(int_map_req_v[650]));
	MUX21X1 U651(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[10]) ,.Q(int_map_req_v[651]));
	MUX21X1 U652(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[10]) ,.Q(int_map_req_v[652]));
	MUX21X1 U653(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[10]) ,.Q(int_map_req_v[653]));
	MUX21X1 U654(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[10]) ,.Q(int_map_req_v[654]));
	MUX21X1 U655(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[10]) ,.Q(int_map_req_v[655]));
	MUX21X1 U656(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[10]) ,.Q(int_map_req_v[656]));
	MUX21X1 U657(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[10]) ,.Q(int_map_req_v[657]));
	MUX21X1 U658(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[10]) ,.Q(int_map_req_v[658]));
	MUX21X1 U659(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[10]) ,.Q(int_map_req_v[659]));
	MUX21X1 U660(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[10]) ,.Q(int_map_req_v[660]));
	MUX21X1 U661(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[10]) ,.Q(int_map_req_v[661]));
	MUX21X1 U662(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[10]) ,.Q(int_map_req_v[662]));
	MUX21X1 U663(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[10]) ,.Q(int_map_req_v[663]));
	MUX21X1 U664(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[10]) ,.Q(int_map_req_v[664]));
	MUX21X1 U665(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[10]) ,.Q(int_map_req_v[665]));
	MUX21X1 U666(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[5]) ,.Q(int_map_req_v[666]));
	MUX21X1 U667(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[5]) ,.Q(int_map_req_v[667]));
	MUX21X1 U668(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[5]) ,.Q(int_map_req_v[668]));
	MUX21X1 U669(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[5]) ,.Q(int_map_req_v[669]));
	MUX21X1 U670(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[5]) ,.Q(int_map_req_v[670]));
	MUX21X1 U671(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[5]) ,.Q(int_map_req_v[671]));
	MUX21X1 U672(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[5]) ,.Q(int_map_req_v[672]));
	MUX21X1 U673(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[5]) ,.Q(int_map_req_v[673]));
	MUX21X1 U674(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[5]) ,.Q(int_map_req_v[674]));
	MUX21X1 U675(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[5]) ,.Q(int_map_req_v[675]));
	MUX21X1 U676(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[5]) ,.Q(int_map_req_v[676]));
	MUX21X1 U677(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[5]) ,.Q(int_map_req_v[677]));
	MUX21X1 U678(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[5]) ,.Q(int_map_req_v[678]));
	MUX21X1 U679(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[5]) ,.Q(int_map_req_v[679]));
	MUX21X1 U680(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[5]) ,.Q(int_map_req_v[680]));
	MUX21X1 U681(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[5]) ,.Q(int_map_req_v[681]));
	MUX21X1 U682(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[5]) ,.Q(int_map_req_v[682]));
	MUX21X1 U683(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[5]) ,.Q(int_map_req_v[683]));
	MUX21X1 U684(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[5]) ,.Q(int_map_req_v[684]));
	MUX21X1 U685(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[5]) ,.Q(int_map_req_v[685]));
	MUX21X1 U686(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[5]) ,.Q(int_map_req_v[686]));
	MUX21X1 U687(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[5]) ,.Q(int_map_req_v[687]));
	MUX21X1 U688(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[5]) ,.Q(int_map_req_v[688]));
	MUX21X1 U689(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[5]) ,.Q(int_map_req_v[689]));
	MUX21X1 U690(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[5]) ,.Q(int_map_req_v[690]));
	MUX21X1 U691(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[5]) ,.Q(int_map_req_v[691]));
	MUX21X1 U692(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[5]) ,.Q(int_map_req_v[692]));
	MUX21X1 U693(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[5]) ,.Q(int_map_req_v[693]));
	MUX21X1 U694(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[5]) ,.Q(int_map_req_v[694]));
	MUX21X1 U695(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[5]) ,.Q(int_map_req_v[695]));
	MUX21X1 U696(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[5]) ,.Q(int_map_req_v[696]));
	MUX21X1 U697(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[5]) ,.Q(int_map_req_v[697]));
	MUX21X1 U698(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[5]) ,.Q(int_map_req_v[698]));
	MUX21X1 U699(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[5]) ,.Q(int_map_req_v[699]));
	MUX21X1 U700(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[5]) ,.Q(int_map_req_v[700]));
	MUX21X1 U701(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[5]) ,.Q(int_map_req_v[701]));
	MUX21X1 U702(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[5]) ,.Q(int_map_req_v[702]));
	MUX21X1 U703(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[0]) ,.Q(int_map_req_v[703]));
	MUX21X1 U704(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[0]) ,.Q(int_map_req_v[704]));
	MUX21X1 U705(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[0]) ,.Q(int_map_req_v[705]));
	MUX21X1 U706(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[0]) ,.Q(int_map_req_v[706]));
	MUX21X1 U707(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[0]) ,.Q(int_map_req_v[707]));
	MUX21X1 U708(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[0]) ,.Q(int_map_req_v[708]));
	MUX21X1 U709(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[0]) ,.Q(int_map_req_v[709]));
	MUX21X1 U710(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[0]) ,.Q(int_map_req_v[710]));
	MUX21X1 U711(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[0]) ,.Q(int_map_req_v[711]));
	MUX21X1 U712(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[0]) ,.Q(int_map_req_v[712]));
	MUX21X1 U713(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[0]) ,.Q(int_map_req_v[713]));
	MUX21X1 U714(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[0]) ,.Q(int_map_req_v[714]));
	MUX21X1 U715(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[0]) ,.Q(int_map_req_v[715]));
	MUX21X1 U716(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[0]) ,.Q(int_map_req_v[716]));
	MUX21X1 U717(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[0]) ,.Q(int_map_req_v[717]));
	MUX21X1 U718(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[0]) ,.Q(int_map_req_v[718]));
	MUX21X1 U719(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[0]) ,.Q(int_map_req_v[719]));
	MUX21X1 U720(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[0]) ,.Q(int_map_req_v[720]));
	MUX21X1 U721(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[0]) ,.Q(int_map_req_v[721]));
	MUX21X1 U722(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[0]) ,.Q(int_map_req_v[722]));
	MUX21X1 U723(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[0]) ,.Q(int_map_req_v[723]));
	MUX21X1 U724(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[0]) ,.Q(int_map_req_v[724]));
	MUX21X1 U725(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[0]) ,.Q(int_map_req_v[725]));
	MUX21X1 U726(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[0]) ,.Q(int_map_req_v[726]));
	MUX21X1 U727(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[0]) ,.Q(int_map_req_v[727]));
	MUX21X1 U728(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[0]) ,.Q(int_map_req_v[728]));
	MUX21X1 U729(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[0]) ,.Q(int_map_req_v[729]));
	MUX21X1 U730(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[0]) ,.Q(int_map_req_v[730]));
	MUX21X1 U731(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[0]) ,.Q(int_map_req_v[731]));
	MUX21X1 U732(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[0]) ,.Q(int_map_req_v[732]));
	MUX21X1 U733(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[0]) ,.Q(int_map_req_v[733]));
	MUX21X1 U734(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[0]) ,.Q(int_map_req_v[734]));
	MUX21X1 U735(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[0]) ,.Q(int_map_req_v[735]));
	MUX21X1 U736(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[0]) ,.Q(int_map_req_v[736]));
	MUX21X1 U737(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[0]) ,.Q(int_map_req_v[737]));
	MUX21X1 U738(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[0]) ,.Q(int_map_req_v[738]));
	MUX21X1 U739(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[0]) ,.Q(int_map_req_v[739]));
	MUX21X1 U33(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[19]), .S(int_route_v[0]) ,.Q(int_resp_v[0]));
	MUX21X1 U34(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[20]), .S(int_route_v[0]) ,.Q(int_resp_v[1]));
	MUX21X1 U35(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[18]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));
	MUX21X1 U36(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[19]), .S(int_route_v[5]) ,.Q(int_resp_v[2]));
	MUX21X1 U37(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[17]), .S(int_route_v[10]) ,.Q(int_resp_v[2]));
	MUX21X1 U38(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[18]), .S(int_route_v[10]) ,.Q(int_resp_v[3]));
	MUX21X1 U39(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[16]), .S(int_route_v[15]) ,.Q(int_resp_v[3]));
	MUX21X1 U40(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[17]), .S(int_route_v[15]) ,.Q(int_resp_v[4]));
	
endmodule 