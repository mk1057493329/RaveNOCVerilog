module router_ravenoc (clk,arst,north_send,north_recv,south_send,south_recv,west_send,west_recv,east_send,east_recv,local_send,local_recv);

	input clk;
	input arst;
	input north_send;
	input west_recv;
	input east_send;
	input east_recv;
	input north_recv;
	input south_send;
	input south_recv;
	input west_send;
	input local_send;
	input local_recv;
	
	wire south_recv_resp,south_recv_req,south_send_resp,south_send_req,west_recv_resp,west_recv_req,west_send_resp,west_send_req,north_recv_resp,north_recv_req,north_send_resp,north_send_req,east_recv_resp,east_recv_req,east_send_resp,east_send_req,local_recv_resp,local_recv_req,local_send_resp,local_send_req;
	wire [194:0] int_req_v;
	wire [4:0] int_resp_v;
	wire [24:0] int_route_v;
	wire [739:0] int_map_req_v;
	wire [19:0] int_map_resp_v;
	wire [194:0] ext_req_v_i;
	wire [4:0] ext_resp_v_o;
	wire [194:0] ext_req_v_o;
	wire [4:0] ext_resp_v_i;
	wire [11:0] valid_from_im_output_module;
	wire [11:0] grant_im_output_module;
	wire [2:0] tail_flit_im_output_module;
	wire [1:0] vc_ch_act_out_output_module;
	wire req_out_output_module,xnor1resu1_output_module,xnor2resu1_output_module,and1resu1_output_module,xor1resu1_output_module,and2resu1_output_module,head_flit_output_module_32_not_output_module,and3resu1_output_module,nor23resu1_output_module,nor23resu2_output_module,and4resu1_output_module,and5resu1_output_module,or12resu12_output_module,nor23resu3_output_module,and6resu1_output_module,nand1resu_output_module,and8resu1_output_module,norfinresu1_output_module,and9resu1_output_module,and10resu1_output_module,and11resu1_output_module;
	wire [33:0] head_flit_output_module;
	wire [1:0] _sv2v_jump_output_module;
	wire [31:0] in_mod_output_module;
	wire [31:0] vc_channel_output_module;
	wire [1:0] _sv2v_jump_output_module_1;
	wire [31:0] i_output_module;
    wire [1:0] mask_ff_rr_arbiter, next_mask_rr_arbiter, mask_req_rr_arbiter, _sv2v_jump_rr_rr_arbiter, i_rr_arbiter, j_rr_arbiter, raw_grant_rr_arbiter, masked_grant_rr_arbiter, temp_mask_ff_rr_arbiter, _sv2v_jump_high_prior_arbiter1, i_high_prior_arbiter1, _sv2v_jump_high_prior_arbiter2, i_high_prior_arbiter2, mask_ff_rr_arbiter1, next_mask_rr_arbiter1, mask_req_rr_arbiter1, _sv2v_jump_rr_rr_arbiter1, i_rr_arbiter1, j_rr_arbiter1, raw_grant_rr_arbiter1, masked_grant_rr_arbiter1, temp_mask_ff_rr_arbiter11, _sv2v_jump_high_prior_arbiter11, i_high_prior_arbiter11, _sv2v_jump_high_prior_arbiter21, i_high_prior_arbiter21,mask_ff_rr_arbiter2,next_mask_rr_arbiter2,mask_req_rr_arbiter2,_sv2v_jump_rr_rr_arbiter2,i_rr_arbiter2,j_rr_arbiter2,raw_grant_rr_arbiter2,masked_grant_rr_arbiter2,temp_mask_ff_rr_arbiter22,_sv2v_jump_high_prior_arbiter12,i_high_prior_arbiter12,_sv2v_jump_high_prior_arbiter22,i_high_prior_arbiter22;

    wire xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter,xnor1res_rr_arbiter,firstif_rr_arbiter,secondif_rr_arbiter,thirdif_rr_arbiter,fourthif_rr_arbiter,not_i_rr_arbiter,arst_value_rr_arbiter,xnores_high_prior_arbiter1,i_0_not_high_prior_arbiter1,nandres_high_prior_arbiter1,xnores_high_prior_arbiter2,i_0_not_high_prior_arbiter2,nandres_high_prior_arbiter2,xnor0res_rr_arbiter1,xnor1res_rr_arbiter1,firstif_rr_arbiter1,secondif_rr_arbiter1,thirdif_rr_arbiter1,fourthif_rr_arbiter1,not_i_rr_arbiter11,arst_value_rr_arbiter1,xnores_high_prior_arbiter11,i_0_not_high_prior_arbiter11,nandres_high_prior_arbiter11,xnores_high_prior_arbiter22,i_0_not_high_prior_arbiter22,nandres_high_prior_arbiter22,xnor0res_rr_arbiter2,xnor1res_rr_arbiter2,firstif_rr_arbiter2,secondif_rr_arbiter2,thirdif_rr_arbiter2,fourthif_rr_arbiter2,not_i_rr_arbiter22,arst_value_rr_arbiter2,xnores_high_prior_arbiter12,i_0_not_high_prior_arbiter12,nandres_high_prior_arbiter12;

    wire [11:0] valid_from_im_output_module1;
    wire [11:0] grant_im_output_module1;
    wire [2:0] tail_flit_im_output_module1;
    wire [1:0] vc_ch_act_out_output_module1;
    wire req_out_output_module1,xnor1resu1_output_module1,xnor2resu1_output_module1,and1resu1_output_module1,xor1resu1_output_module1,and2resu1_output_module1,head_flit_output_module1_32_not_output_module1,and3resu1_output_module1,nor23resu1_output_module1,nor23resu2_output_module1,and4resu1_output_module1,and5resu1_output_module1,or12resu12_output_module1,nor23resu3_output_module1,and6resu1_output_module1,nand1resu_output_module1,and8resu1_output_module1,norfinresu1_output_module1,and9resu1_output_module1,and10resu1_output_module1,and11resu1_output_module1;
    wire [33:0] head_flit_output_module1;
    wire [1:0] _sv2v_jump_output_module1;
    wire [31:0] in_mod_output_module1;
    wire [31:0] vc_channel_output_module1;
    wire [1:0] _sv2v_jump_output_module1_1;
    wire [31:0] i_output_module1;
    wire [1:0] mask_ff_rr_arbiter11, next_mask_rr_arbiter11, mask_req_rr_arbiter11, _sv2v_jump_rr_rr_arbiter11, i_rr_arbiter11, j_rr_arbiter11, raw_grant_rr_arbiter11, masked_grant_rr_arbiter11, temp_mask_ff_rr_arbiter1111, _sv2v_jump_high_prior_arbiter111, i_high_prior_arbiter111, _sv2v_jump_high_prior_arbiter211, i_high_prior_arbiter211, mask_ff_rr_arbiter111, next_mask_rr_arbiter111, mask_req_rr_arbiter111, _sv2v_jump_rr_rr_arbiter111, i_rr_arbiter111, j_rr_arbiter111, raw_grant_rr_arbiter111, masked_grant_rr_arbiter111, temp_mask_ff_rr_arbiter111111, _sv2v_jump_high_prior_arbiter1111, i_high_prior_arbiter1111, _sv2v_jump_high_prior_arbiter2111, i_high_prior_arbiter2111,mask_ff_rr_arbiter112,next_mask_rr_arbiter112,mask_req_rr_arbiter112,_sv2v_jump_rr_rr_arbiter112,i_rr_arbiter112,j_rr_arbiter112,raw_grant_rr_arbiter112,masked_grant_rr_arbiter112,temp_mask_ff_rr_arbiter111122,_sv2v_jump_high_prior_arbiter1112,i_high_prior_arbiter1112,_sv2v_jump_high_prior_arbiter2112,i_high_prior_arbiter2112;

    wire xnores_high_prior_arbiter2111,i_0_not_high_prior_arbiter2111,nandres_high_prior_arbiter2111,xnor0res_rr_arbiter11,xnor1res_rr_arbiter11,firstif_rr_arbiter11,secondif_rr_arbiter11,thirdif_rr_arbiter11,fourthif_rr_arbiter11,not_i_rr_arbiter1111,arst_value_rr_arbiter11,xnores_high_prior_arbiter111,i_0_not_high_prior_arbiter111,nandres_high_prior_arbiter111,xnores_high_prior_arbiter21,i_0_not_high_prior_arbiter21,nandres_high_prior_arbiter21,xnor0res_rr_arbiter111,xnor1res_rr_arbiter111,firstif_rr_arbiter111,secondif_rr_arbiter111,thirdif_rr_arbiter111,fourthif_rr_arbiter111,not_i_rr_arbiter111111,arst_value_rr_arbiter111,xnores_high_prior_arbiter1111,i_0_not_high_prior_arbiter1111,nandres_high_prior_arbiter1111,xnores_high_prior_arbiter212,i_0_not_high_prior_arbiter212,nandres_high_prior_arbiter212,xnor0res_rr_arbiter112,xnor1res_rr_arbiter112,firstif_rr_arbiter112,secondif_rr_arbiter112,thirdif_rr_arbiter112,fourthif_rr_arbiter112,not_i_rr_arbiter111122,arst_value_rr_arbiter112,xnores_high_prior_arbiter1112,i_0_not_high_prior_arbiter1112,nandres_high_prior_arbiter1112;

    wire [11:0] valid_from_im_output_module2;
    wire [11:0] grant_im_output_module2;
    wire [2:0] tail_flit_im_output_module2;
    wire [1:0] vc_ch_act_out_output_module2;
    wire req_out_output_module2,xnor1resu1_output_module2,xnor2resu1_output_module2,and1resu1_output_module2,xor1resu1_output_module2,and2resu1_output_module2,head_flit_output_module2_32_not_output_module2,and3resu1_output_module2,nor23resu1_output_module2,nor23resu2_output_module2,and4resu1_output_module2,and5resu1_output_module2,or12resu12_output_module2,nor23resu3_output_module2,and6resu1_output_module2,nand1resu_output_module2,and8resu1_output_module2,norfinresu1_output_module2,and9resu1_output_module2,and10resu1_output_module2,and11resu1_output_module2;
    wire [33:0] head_flit_output_module2;
    wire [1:0] _sv2v_jump_output_module2;
    wire [31:0] in_mod_output_module2;
    wire [31:0] vc_channel_output_module2;
    wire [1:0] _sv2v_jump_output_module2_1;
    wire [31:0] i_output_module2;
    wire [1:0] mask_ff_rr_arbiter22, next_mask_rr_arbiter22, mask_req_rr_arbiter22, _sv2v_jump_rr_rr_arbiter22, i_rr_arbiter22, j_rr_arbiter22, raw_grant_rr_arbiter22, masked_grant_rr_arbiter22, temp_mask_ff_rr_arbiter2222, _sv2v_jump_high_prior_arbiter122, i_high_prior_arbiter122, _sv2v_jump_high_prior_arbiter222, i_high_prior_arbiter222, mask_ff_rr_arbiter221, next_mask_rr_arbiter221, mask_req_rr_arbiter221, _sv2v_jump_rr_rr_arbiter221, i_rr_arbiter221, j_rr_arbiter221, raw_grant_rr_arbiter221, masked_grant_rr_arbiter221, temp_mask_ff_rr_arbiter222211, _sv2v_jump_high_prior_arbiter1221, i_high_prior_arbiter1221, _sv2v_jump_high_prior_arbiter2221, i_high_prior_arbiter2221,mask_ff_rr_arbiter222,next_mask_rr_arbiter222,mask_req_rr_arbiter222,_sv2v_jump_rr_rr_arbiter222,i_rr_arbiter222,j_rr_arbiter222,raw_grant_rr_arbiter222,masked_grant_rr_arbiter222,temp_mask_ff_rr_arbiter222222,_sv2v_jump_high_prior_arbiter1222,i_high_prior_arbiter1222,_sv2v_jump_high_prior_arbiter2222,i_high_prior_arbiter2222;

    wire xnores_high_prior_arbiter22212,i_0_not_high_prior_arbiter22212,nandres_high_prior_arbiter22212,xnor0res_rr_arbiter22,xnor1res_rr_arbiter22,firstif_rr_arbiter22,secondif_rr_arbiter22,thirdif_rr_arbiter22,fourthif_rr_arbiter22,not_i_rr_arbiter2222,arst_value_rr_arbiter22,xnores_high_prior_arbiter122,i_0_not_high_prior_arbiter122,nandres_high_prior_arbiter122,xnores_high_prior_arbiter222,i_0_not_high_prior_arbiter222,nandres_high_prior_arbiter222,xnor0res_rr_arbiter221,xnor1res_rr_arbiter221,firstif_rr_arbiter221,secondif_rr_arbiter221,thirdif_rr_arbiter221,fourthif_rr_arbiter221,not_i_rr_arbiter222211,arst_value_rr_arbiter221,xnores_high_prior_arbiter1221,i_0_not_high_prior_arbiter1221,nandres_high_prior_arbiter1221,xnores_high_prior_arbiter2222,i_0_not_high_prior_arbiter2222,nandres_high_prior_arbiter2222,xnor0res_rr_arbiter222,xnor1res_rr_arbiter222,firstif_rr_arbiter222,secondif_rr_arbiter222,thirdif_rr_arbiter222,fourthif_rr_arbiter222,not_i_rr_arbiter222222,arst_value_rr_arbiter222,xnores_high_prior_arbiter1222,i_0_not_high_prior_arbiter1222,nandres_high_prior_arbiter1222;


    wire [11:0] valid_from_im_output_module3;
    wire [11:0] grant_im_output_module3;
    wire [2:0] tail_flit_im_output_module3;
    wire [1:0] vc_ch_act_out_output_module3;
    wire req_out_output_module3,xnor1resu1_output_module3,xnor2resu1_output_module3,and1resu1_output_module3,xor1resu1_output_module3,and2resu1_output_module3,head_flit_output_module3_32_not_output_module3,and3resu1_output_module3,nor23resu1_output_module3,nor23resu2_output_module3,and4resu1_output_module3,and5resu1_output_module3,or12resu12_output_module3,nor23resu3_output_module3,and6resu1_output_module3,nand1resu_output_module3,and8resu1_output_module3,norfinresu1_output_module3,and9resu1_output_module3,and10resu1_output_module3,and11resu1_output_module3;
    wire [33:0] head_flit_output_module3;
    wire [1:0] _sv2v_jump_output_module3;
    wire [31:0] in_mod_output_module3;
    wire [31:0] vc_channel_output_module3;
    wire [1:0] _sv2v_jump_output_module3_1;
    wire [31:0] i_output_module3;
    wire [1:0] mask_ff_rr_arbiter3, next_mask_rr_arbiter3, mask_req_rr_arbiter3, _sv2v_jump_rr_rr_arbiter3, i_rr_arbiter3, j_rr_arbiter3, raw_grant_rr_arbiter3, masked_grant_rr_arbiter3, temp_mask_ff_rr_arbiter33, _sv2v_jump_high_prior_arbiter13, i_high_prior_arbiter13, _sv2v_jump_high_prior_arbiter23, i_high_prior_arbiter23, mask_ff_rr_arbiter31, next_mask_rr_arbiter31, mask_req_rr_arbiter31, _sv2v_jump_rr_rr_arbiter31, i_rr_arbiter31, j_rr_arbiter31, raw_grant_rr_arbiter31, masked_grant_rr_arbiter31, temp_mask_ff_rr_arbiter3311, _sv2v_jump_high_prior_arbiter131, i_high_prior_arbiter131, _sv2v_jump_high_prior_arbiter231, i_high_prior_arbiter231,mask_ff_rr_arbiter32,next_mask_rr_arbiter32,mask_req_rr_arbiter32,_sv2v_jump_rr_rr_arbiter32,i_rr_arbiter32,j_rr_arbiter32,raw_grant_rr_arbiter32,masked_grant_rr_arbiter32,temp_mask_ff_rr_arbiter3322,_sv2v_jump_high_prior_arbiter132,i_high_prior_arbiter132,_sv2v_jump_high_prior_arbiter232,i_high_prior_arbiter232;

    wire xnores_high_prior_arbiter2313,i_0_not_high_prior_arbiter2313,nandres_high_prior_arbiter2313,xnor0res_rr_arbiter3,xnor1res_rr_arbiter3,firstif_rr_arbiter3,secondif_rr_arbiter3,thirdif_rr_arbiter3,fourthif_rr_arbiter3,not_i_rr_arbiter33,arst_value_rr_arbiter3,xnores_high_prior_arbiter13,i_0_not_high_prior_arbiter13,nandres_high_prior_arbiter13,xnores_high_prior_arbiter23,i_0_not_high_prior_arbiter23,nandres_high_prior_arbiter23,xnor0res_rr_arbiter31,xnor1res_rr_arbiter31,firstif_rr_arbiter31,secondif_rr_arbiter31,thirdif_rr_arbiter31,fourthif_rr_arbiter31,not_i_rr_arbiter3311,arst_value_rr_arbiter31,xnores_high_prior_arbiter131,i_0_not_high_prior_arbiter131,nandres_high_prior_arbiter131,xnores_high_prior_arbiter232,i_0_not_high_prior_arbiter232,nandres_high_prior_arbiter232,xnor0res_rr_arbiter32,xnor1res_rr_arbiter32,firstif_rr_arbiter32,secondif_rr_arbiter32,thirdif_rr_arbiter32,fourthif_rr_arbiter32,not_i_rr_arbiter3322,arst_value_rr_arbiter32,xnores_high_prior_arbiter132,i_0_not_high_prior_arbiter132,nandres_high_prior_arbiter132;


    wire [11:0] valid_from_im_output_module4;
    wire [11:0] grant_im_output_module4;
    wire [2:0] tail_flit_im_output_module4;
    wire [1:0] vc_ch_act_out_output_module4;
    wire req_out_output_module4,xnor1resu1_output_module4,xnor2resu1_output_module4,and1resu1_output_module4,xor1resu1_output_module4,and2resu1_output_module4,head_flit_output_module4_32_not_output_module4,and3resu1_output_module4,nor23resu1_output_module4,nor23resu2_output_module4,and4resu1_output_module4,and5resu1_output_module4,or12resu12_output_module4,nor23resu3_output_module4,and6resu1_output_module4,nand1resu_output_module4,and8resu1_output_module4,norfinresu1_output_module4,and9resu1_output_module4,and10resu1_output_module4,and11resu1_output_module4;
    wire [33:0] head_flit_output_module4;
    wire [1:0] _sv2v_jump_output_module4;
    wire [31:0] in_mod_output_module4;
    wire [31:0] vc_channel_output_module4;
    wire [1:0] _sv2v_jump_output_module4_1;
    wire [31:0] i_output_module4;
    wire [1:0] mask_ff_rr_arbiter4, next_mask_rr_arbiter4, mask_req_rr_arbiter4, _sv2v_jump_rr_rr_arbiter4, i_rr_arbiter4, j_rr_arbiter4, raw_grant_rr_arbiter4, masked_grant_rr_arbiter4, temp_mask_ff_rr_arbiter44, _sv2v_jump_high_prior_arbiter14, i_high_prior_arbiter14, _sv2v_jump_high_prior_arbiter24, i_high_prior_arbiter24, mask_ff_rr_arbiter41, next_mask_rr_arbiter41, mask_req_rr_arbiter41, _sv2v_jump_rr_rr_arbiter41, i_rr_arbiter41, j_rr_arbiter41, raw_grant_rr_arbiter41, masked_grant_rr_arbiter41, temp_mask_ff_rr_arbiter4411, _sv2v_jump_high_prior_arbiter141, i_high_prior_arbiter141, _sv2v_jump_high_prior_arbiter241, i_high_prior_arbiter241,mask_ff_rr_arbiter42,next_mask_rr_arbiter42,mask_req_rr_arbiter42,_sv2v_jump_rr_rr_arbiter42,i_rr_arbiter42,j_rr_arbiter42,raw_grant_rr_arbiter42,masked_grant_rr_arbiter42,temp_mask_ff_rr_arbiter4422,_sv2v_jump_high_prior_arbiter142,i_high_prior_arbiter142,_sv2v_jump_high_prior_arbiter242,i_high_prior_arbiter242;

    wire xnores_high_prior_arbiter2414,i_0_not_high_prior_arbiter2414,nandres_high_prior_arbiter2414,xnor0res_rr_arbiter4,xnor1res_rr_arbiter4,firstif_rr_arbiter4,secondif_rr_arbiter4,thirdif_rr_arbiter4,fourthif_rr_arbiter4,not_i_rr_arbiter44,arst_value_rr_arbiter4,xnores_high_prior_arbiter14,i_0_not_high_prior_arbiter14,nandres_high_prior_arbiter14,xnores_high_prior_arbiter24,i_0_not_high_prior_arbiter24,nandres_high_prior_arbiter24,xnor0res_rr_arbiter41,xnor1res_rr_arbiter41,firstif_rr_arbiter41,secondif_rr_arbiter41,thirdif_rr_arbiter41,fourthif_rr_arbiter41,not_i_rr_arbiter4411,arst_value_rr_arbiter41,xnores_high_prior_arbiter141,i_0_not_high_prior_arbiter141,nandres_high_prior_arbiter141,xnores_high_prior_arbiter242,i_0_not_high_prior_arbiter242,nandres_high_prior_arbiter242,xnor0res_rr_arbiter42,xnor1res_rr_arbiter42,firstif_rr_arbiter42,secondif_rr_arbiter42,thirdif_rr_arbiter42,fourthif_rr_arbiter42,not_i_rr_arbiter4422,arst_value_rr_arbiter42,xnores_high_prior_arbiter142,i_0_not_high_prior_arbiter142,nandres_high_prior_arbiter142;

   	wire [8:0] routing_table_ff_input_router;
	wire [2:0] next_rt_input_router;
	wire [33:0] flit_input_router;
	wire new_rt_input_router,new_rt_input_routernot,norres_1_input_router,norres_2_input_router,norres_3_input_router,andfinres_input_router,and2result_input_router,norres_4_input_router,invres1_input_router,invres2_input_router,and3result_input_router,and4result_input_router,and5result_input_router,norres_5_input_router,and6result_input_router,and7result_input_router,and8result_input_router,and9result_input_router,and10result_input_router,and11result_input_router,orres1_input_router,orres2_input_router,orres3_input_router,finand1_input_router,finand2_input_router,finand3_input_router,nextrt2not_input_router,secondAndc_input_router,norres_5_input_router_2,and62result_input_router,and7result_input_router2,orres1_input_router2,finand1_input_router2,finand2_input_router2,and8result_input_router2,orres2_input_router2,and9result_input_router2,orres3_input_router2,finand3_input_router2,and11result_input_router2,nextrt2not_input_router,and10result_input_router2,arst_valuenot_input_router,finand3_input_router22;
    
    wire [8:0] routing_table_ff_input_router1;
    wire [2:0] next_rt_input_router1;
    wire [33:0] flit_input_router1;
    wire new_rt_input_router1,new_rt_input_router1not,norres_1_input_router1,norres_2_input_router1,norres_3_input_router1,andfinres_input_router1,and2result_input_router1,norres_4_input_router1,invres1_input_router1,invres2_input_router1,and3result_input_router1,and4result_input_router1,and5result_input_router1,norres_5_input_router1,and6result_input_router1,and7result_input_router1,and8result_input_router1,and9result_input_router1,and10result_input_router1,and11result_input_router1,orres1_input_router1,orres2_input_router1,orres3_input_router1,finand1_input_router1,finand2_input_router1,finand3_input_router1,nextrt2not_input_router11,secondAndc_input_router1,norres_5_input_router1_2,and62result_input_router1,and7result_input_router12,orres1_input_router12,finand1_input_router12,finand2_input_router12,and8result_input_router12,orres2_input_router12,and9result_input_router12,orres3_input_router12,finand3_input_router12,and11result_input_router12,nextrt2not_input_router11,and10result_input_router12,arst_valuenot_input_router1,finand3_input_router122;


    wire [8:0] routing_table_ff_input_router2;
    wire [2:0] next_rt_input_router2;
    wire [33:0] flit_input_router2;
    wire new_rt_input_router2,new_rt_input_router2not,norres_1_input_router2,norres_2_input_router2,norres_3_input_router2,andfinres_input_router2,and2result_input_router2,norres_4_input_router2,invres1_input_router2,invres2_input_router2,and3result_input_router2,and4result_input_router2,and5result_input_router2,norres_5_input_router2,and6result_input_router2,and7result_input_router22,and8result_input_router22,and9result_input_router22,and10result_input_router22,and11result_input_router22,orres1_input_router22,orres2_input_router22,orres3_input_router22,finand1_input_router22,finand2_input_router22,finand3_input_router222,nextrt2not_input_router22,secondAndc_input_router2,norres_5_input_router2_2,and62result_input_router2,and7result_input_router222,orres1_input_router222,finand1_input_router222,finand2_input_router222,and8result_input_router222,orres2_input_router222,and9result_input_router222,orres3_input_router222,finand3_input_router2222,and11result_input_router222,nextrt2not_input_router22,and10result_input_router222,arst_valuenot_input_router2,finand3_input_router22222;


    wire [8:0] routing_table_ff_input_router3;
    wire [2:0] next_rt_input_router3;
    wire [33:0] flit_input_router3;
    wire new_rt_input_router3,new_rt_input_router3not,norres_1_input_router3,norres_2_input_router3,norres_3_input_router3,andfinres_input_router3,and2result_input_router3,norres_4_input_router3,invres1_input_router3,invres2_input_router3,and3result_input_router3,and4result_input_router3,and5result_input_router3,norres_5_input_router3,and6result_input_router3,and7result_input_router3,and8result_input_router3,and9result_input_router3,and10result_input_router3,and11result_input_router3,orres1_input_router3,orres2_input_router3,orres3_input_router3,finand1_input_router3,finand2_input_router3,finand3_input_router3,nextrt2not_input_router33,secondAndc_input_router3,norres_5_input_router3_2,and62result_input_router3,and7result_input_router32,orres1_input_router32,finand1_input_router32,finand2_input_router32,and8result_input_router32,orres2_input_router32,and9result_input_router32,orres3_input_router32,finand3_input_router32,and11result_input_router32,nextrt2not_input_router33,and10result_input_router32,arst_valuenot_input_router3,finand3_input_router322;


    wire [8:0] routing_table_ff_input_router4;
    wire [2:0] next_rt_input_router4;
    wire [33:0] flit_input_router4;
    wire new_rt_input_router4,new_rt_input_router4not,norres_1_input_router4,norres_2_input_router4,norres_3_input_router4,andfinres_input_router4,and2result_input_router4,norres_4_input_router4,invres1_input_router4,invres2_input_router4,and3result_input_router4,and4result_input_router4,and5result_input_router4,norres_5_input_router4,and6result_input_router4,and7result_input_router4,and8result_input_router4,and9result_input_router4,and10result_input_router4,and11result_input_router4,orres1_input_router4,orres2_input_router4,orres3_input_router4,finand1_input_router4,finand2_input_router4,finand3_input_router4,nextrt2not_input_router44,secondAndc_input_router4,norres_5_input_router4_2,and62result_input_router4,and7result_input_router42,orres1_input_router42,finand1_input_router42,finand2_input_router42,and8result_input_router42,orres2_input_router42,and9result_input_router42,orres3_input_router42,finand3_input_router42,and11result_input_router42,nextrt2not_input_router44,and10result_input_router42,arst_valuenot_input_router4,finand3_input_router422;

	wire [110:0] from_input_req_in_jump_input_datapathput_datapath;
	wire [2:0] from_input_resp_input_datapath;
	wire [110:0] to_output_req_in_jump_input_datapathput_datapath;
	wire [2:0] to_output_resp_input_datapath;
	wire [1:0] vc_ch_act_in_input_datapath;
	wire [1:0] vc_ch_act_out_input_datapath;
	wire [2:0] i_input_datapath;
	wire [2:0] j_input_datapath;
	wire [0:1] _sv2v_jump_input_datapath;

	wire req_in_jump_input_datapath,req_out_jump_input_datapath,xnor1resu_input_datapath,xnor2resu_input_datapath,and1resu_input_datapath,cond1line_input_datapath,req_in_jump_input_datapath_not,and2resu_input_datapath,xor1resu_input_datapath,nand1resu_input_datapath,xnor23resu_input_datapath,and4resu_input_datapath,write_flit_vc_buffer,norres_vc_buffer_vc_buffer,full_vc_buffer,empty_vc_buffer,error_vc_buffer,read_flit_vc_buffer,locked_by_route_ff_vc_buffer,next_locked_vc_buffer,orres_vc_buffer,or1res_vc_buffer,or2res_vc_buffer,finres1_vc_buffer,andres1_vc_buffer,full_vc_buffer_not,locked_by_route_ff_vc_buffer_not,thirdand_vc_buffer,u1temp_fifomodule,u2temp_fifomodule,u4temp_fifomodule,full_vc_buffer_not_fifomodule,u7temp_fifomodule,u9temp_fifomodule,u10carry_fifomodule,u11carry_fifomodule,empty_vc_buffer_not_fifomodule,u13temp_fifomodule,u14temp_fifomodule,u15carry_fifomodule,u16carry_fifomodule,u17res_fifomodule,u18res_fifomodule,write_ptr_ff_fifomodule_0_not,write_ptr_ff_fifomodule_1_not,b0wire_fifomodule,b1wire_fifomodule,u23temp_fifomodule_not_fifomodule,u23temp_fifomodule,boutb_fifomodule,bouta_fifomodule,boutmain_fifomodule,arst_value_fifomodule,write_flit1_vc_buffer1,norres_vc_buffer1_vc_buffer1,full_vc_buffer1,empty_vc_buffer1,error_vc_buffer1,read_flit1_vc_buffer1,locked_by_route_ff_vc_buffer1,next_locked_vc_buffer1,orres_vc_buffer1,or1res_vc_buffer1,or2res_vc_buffer1,finres1_vc_buffer1,andres1_vc_buffer1,full_vc_buffer1_not1,locked_by_route_ff_vc_buffer1_not1,thirdand_vc_buffer1,u1temp_fifomodule1,u2temp_fifomodule1,u4temp_fifomodule1,full_vc_buffer1_not1_fifomodule1,u7temp_fifomodule1,u9temp_fifomodule1,u10carry_fifomodule1,u11carry_fifomodule1,empty_vc_buffer1_not_fifomodule1,u13temp_fifomodule1,u14temp_fifomodule1,u15carry_fifomodule1,u16carry_fifomodule1,u17res_fifomodule1,u18res_fifomodule1,write_ptr_ff_fifomodule1_0_not1,write_ptr_ff_fifomodule1_1_not1,b0wire_fifomodule1,b1wire_fifomodule1,u23temp_fifomodule1_not_fifomodule1,u23temp_fifomodule1,boutb_fifomodule1,bouta_fifomodule1,boutmain_fifomodule1,arst_value_fifomodule1,write_flit2_vc_buffer2,norres_vc_buffer2_vc_buffer2,full_vc_buffer2,empty_vc_buffer2,error_vc_buffer2,read_flit2_vc_buffer2,locked_by_route_ff_vc_buffer2,next_locked_vc_buffer2,orres_vc_buffer2,or1res_vc_buffer2,or2res_vc_buffer2,finres1_vc_buffer2,andres1_vc_buffer2,full_vc_buffer2_not2,locked_by_route_ff_vc_buffer2_not2,thirdand_vc_buffer2,u1temp_fifomodule2,u2temp_fifomodule2,u4temp_fifomodule2,full_vc_buffer2_not2_fifomodule2,u7temp_fifomodule2,u9temp_fifomodule2,u10carry_fifomodule2,u11carry_fifomodule2,empty_vc_buffer2_not_fifomodule2,u13temp_fifomodule2,u14temp_fifomodule2,u15carry_fifomodule2,u16carry_fifomodule2,u17res_fifomodule2,u18res_fifomodule2,write_ptr_ff_fifomodule2_0_not2,write_ptr_ff_fifomodule2_1_not2,b0wire_fifomodule2,b1wire_fifomodule2,u23temp_fifomodule2_not_fifomodule2,u23temp_fifomodule2,boutb_fifomodule2,bouta_fifomodule2,boutmain_fifomodule2,arst_value_fifomodule2;
	wire [33:0] flit,flit1,flit2;
	wire [15:0] fifo_ff_fifomodule,fifo_ff_fifomodule1,fifo_ff_fifomodule2;
	wire [1:0] write_ptr_ff_fifomodule,read_ptr_ff_fifomodule,next_write_ptr_fifomodule,next_read_ptr_fifomodule,fifo_ocup_fifomodule,write_ptr_ff_fifomodule1,read_ptr_ff_fifomodule1,next_write_ptr_fifomodule1,next_read_ptr_fifomodule1,fifo_ocup_fifomodule1,write_ptr_ff_fifomodule2,read_ptr_ff_fifomodule2,next_write_ptr_fifomodule2,next_read_ptr_fifomodule2,fifo_ocup_fifomodule2;

	wire [110:0] from_input_req_in_jump_input_datapath1put_datapath1;
	wire [2:0] from_input_resp_input_datapath1;
	wire [110:0] to_output_req_in_jump_input_datapath1put_datapath1;
	wire [2:0] to_output_resp_input_datapath1;
	wire [1:0] vc_ch_act_in_input_datapath1;
	wire [1:0] vc_ch_act_out_input_datapath1;
	wire [2:0] i_input_datapath1;
	wire [2:0] j_input_datapath1;
	wire [0:1] _sv2v_jump_input_datapath1;

	wire req_in_jump_input_datapath1,req_out_jump_input_datapath1,xnor1resu_input_datapath1,xnor2resu_input_datapath1,and1resu_input_datapath1,cond1line_input_datapath1,req_in_jump_input_datapath1_not,and2resu_input_datapath1,xor1resu_input_datapath1,nand1resu_input_datapath11,xnor23resu_input_datapath1,and4resu_input_datapath1,write_flit11_vc_buffer1,norres_vc_buffer11_vc_buffer11,full_vc_buffer11,empty_vc_buffer11,error_vc_buffer11,read_flit11_vc_buffer1,locked_by_route_ff_vc_buffer11,next_locked_vc_buffer11,orres_vc_buffer11,or1res_vc_buffer11,or2res_vc_buffer11,finres1_vc_buffer11,andres1_vc_buffer11,full_vc_buffer11_not,locked_by_route_ff_vc_buffer11_not,thirdand_vc_buffer11,u1temp_fifomodule11,u2temp_fifomodule11,u4temp_fifomodule11,full_vc_buffer11_not_fifomodule,u7temp_fifomodule11,u9temp_fifomodule11,u10carry_fifomodule11,u11carry_fifomodule11,empty_vc_buffer11_not_fifomodule,u13temp_fifomodule11,u14temp_fifomodule11,u15carry_fifomodule11,u16carry_fifomodule11,u17res_fifomodule11,u18res_fifomodule11,write_ptr_ff_fifomodule11_0_not1,write_ptr_ff_fifomodule11_1_not1,b0wire_fifomodule11,b1wire_fifomodule11,u23temp_fifomodule11_not_fifomodule11,u23temp_fifomodule11,boutb_fifomodule11,bouta_fifomodule11,boutmain_fifomodule11,arst_value_fifomodule11,write_flit111_vc_buffer11,norres_vc_buffer111_vc_buffer1,full_vc_buffer111,empty_vc_buffer111,error_vc_buffer111,read_flit111_vc_buffer11,locked_by_route_ff_vc_buffer111,next_locked_vc_buffer111,orres_vc_buffer111,or1res_vc_buffer111,or2res_vc_buffer111,finres1_vc_buffer111,andres1_vc_buffer111,full_vc_buffer111_not1,locked_by_route_ff_vc_buffer111_not1,thirdand_vc_buffer111,u1temp_fifomodule111,u2temp_fifomodule111,u4temp_fifomodule111,full_vc_buffer111_not1_fifomodule1,u7temp_fifomodule111,u9temp_fifomodule111,u10carry_fifomodule111,u11carry_fifomodule111,empty_vc_buffer111_not_fifomodule1,u13temp_fifomodule111,u14temp_fifomodule111,u15carry_fifomodule111,u16carry_fifomodule111,u17res_fifomodule111,u18res_fifomodule111,write_ptr_ff_fifomodule111_0_not11,write_ptr_ff_fifomodule111_1_not11,b0wire_fifomodule111,b1wire_fifomodule111,u23temp_fifomodule111_not_fifomodule1,u23temp_fifomodule111,boutb_fifomodule111,bouta_fifomodule111,boutmain_fifomodule111,arst_value_fifomodule111,write_flit112_vc_buffer21,norres_vc_buffer112_vc_buffer2,full_vc_buffer112,empty_vc_buffer112,error_vc_buffer112,read_flit112_vc_buffer21,locked_by_route_ff_vc_buffer112,next_locked_vc_buffer112,orres_vc_buffer112,or1res_vc_buffer112,or2res_vc_buffer112,finres1_vc_buffer112,andres1_vc_buffer112,full_vc_buffer112_not2,locked_by_route_ff_vc_buffer112_not2,thirdand_vc_buffer112,u1temp_fifomodule112,u2temp_fifomodule112,u4temp_fifomodule112,full_vc_buffer112_not2_fifomodule2,u7temp_fifomodule112,u9temp_fifomodule112,u10carry_fifomodule112,u11carry_fifomodule112,empty_vc_buffer112_not_fifomodule2,u13temp_fifomodule112,u14temp_fifomodule112,u15carry_fifomodule112,u16carry_fifomodule112,u17res_fifomodule112,u18res_fifomodule112,write_ptr_ff_fifomodule112_0_not21,write_ptr_ff_fifomodule112_1_not21,b0wire_fifomodule112,b1wire_fifomodule112,u23temp_fifomodule112_not_fifomodule2,u23temp_fifomodule112,boutb_fifomodule112,bouta_fifomodule112,boutmain_fifomodule112,arst_value_fifomodule112;
	wire [33:0] flit11,flit111,flit112;
	wire [15:0] fifo_ff_fifomodule11,fifo_ff_fifomodule111,fifo_ff_fifomodule112;
	wire [1:0] write_ptr_ff_fifomodule11,read_ptr_ff_fifomodule11,next_write_ptr_fifomodule11,next_read_ptr_fifomodule11,fifo_ocup_fifomodule11,write_ptr_ff_fifomodule111,read_ptr_ff_fifomodule111,next_write_ptr_fifomodule111,next_read_ptr_fifomodule111,fifo_ocup_fifomodule111,write_ptr_ff_fifomodule112,read_ptr_ff_fifomodule112,next_write_ptr_fifomodule112,next_read_ptr_fifomodule112,fifo_ocup_fifomodule112;

	wire [110:0] from_input_req_in_jump_input_datapath2put_datapath2;
	wire [2:0] from_input_resp_input_datapath2;
	wire [110:0] to_output_req_in_jump_input_datapath2put_datapath2;
	wire [2:0] to_output_resp_input_datapath2;
	wire [1:0] vc_ch_act_in_input_datapath2;
	wire [1:0] vc_ch_act_out_input_datapath2;
	wire [2:0] i_input_datapath2;
	wire [2:0] j_input_datapath2;
	wire [0:1] _sv2v_jump_input_datapath2;

	wire req_in_jump_input_datapath2,req_out_jump_input_datapath2,xnor1resu_input_datapath2,xnor2resu_input_datapath2,and1resu_input_datapath2,cond1line_input_datapath2,req_in_jump_input_datapath2_not,and2resu_input_datapath2,xor1resu_input_datapath2,nand1resu_input_datapath22,xnor23resu_input_datapath2,and4resu_input_datapath2,write_flit22_vc_buffer2,norres_vc_buffer22_vc_buffer22,full_vc_buffer22,empty_vc_buffer22,error_vc_buffer22,read_flit22_vc_buffer2,locked_by_route_ff_vc_buffer22,next_locked_vc_buffer22,orres_vc_buffer22,or1res_vc_buffer22,or2res_vc_buffer22,finres1_vc_buffer22,andres1_vc_buffer22,full_vc_buffer22_not,locked_by_route_ff_vc_buffer22_not,thirdand_vc_buffer22,u1temp_fifomodule22,u2temp_fifomodule22,u4temp_fifomodule22,full_vc_buffer22_not_fifomodule,u7temp_fifomodule22,u9temp_fifomodule22,u10carry_fifomodule22,u11carry_fifomodule22,empty_vc_buffer22_not_fifomodule,u13temp_fifomodule22,u14temp_fifomodule22,u15carry_fifomodule22,u16carry_fifomodule22,u17res_fifomodule22,u18res_fifomodule22,write_ptr_ff_fifomodule22_0_not2,write_ptr_ff_fifomodule22_1_not2,b0wire_fifomodule22,b1wire_fifomodule22,u23temp_fifomodule22_not_fifomodule22,u23temp_fifomodule22,boutb_fifomodule22,bouta_fifomodule22,boutmain_fifomodule22,arst_value_fifomodule22,write_flit221_vc_buffer12,norres_vc_buffer221_vc_buffer1,full_vc_buffer221,empty_vc_buffer221,error_vc_buffer221,read_flit221_vc_buffer12,locked_by_route_ff_vc_buffer221,next_locked_vc_buffer221,orres_vc_buffer221,or1res_vc_buffer221,or2res_vc_buffer221,finres1_vc_buffer221,andres1_vc_buffer221,full_vc_buffer221_not1,locked_by_route_ff_vc_buffer221_not1,thirdand_vc_buffer221,u1temp_fifomodule221,u2temp_fifomodule221,u4temp_fifomodule221,full_vc_buffer221_not1_fifomodule1,u7temp_fifomodule221,u9temp_fifomodule221,u10carry_fifomodule221,u11carry_fifomodule221,empty_vc_buffer221_not_fifomodule1,u13temp_fifomodule221,u14temp_fifomodule221,u15carry_fifomodule221,u16carry_fifomodule221,u17res_fifomodule221,u18res_fifomodule221,write_ptr_ff_fifomodule221_0_not12,write_ptr_ff_fifomodule221_1_not12,b0wire_fifomodule221,b1wire_fifomodule221,u23temp_fifomodule221_not_fifomodule1,u23temp_fifomodule221,boutb_fifomodule221,bouta_fifomodule221,boutmain_fifomodule221,arst_value_fifomodule221,write_flit222_vc_buffer22,norres_vc_buffer222_vc_buffer2,full_vc_buffer222,empty_vc_buffer222,error_vc_buffer222,read_flit222_vc_buffer22,locked_by_route_ff_vc_buffer222,next_locked_vc_buffer222,orres_vc_buffer222,or1res_vc_buffer222,or2res_vc_buffer222,finres1_vc_buffer222,andres1_vc_buffer222,full_vc_buffer222_not2,locked_by_route_ff_vc_buffer222_not2,thirdand_vc_buffer222,u1temp_fifomodule222,u2temp_fifomodule222,u4temp_fifomodule222,full_vc_buffer222_not2_fifomodule2,u7temp_fifomodule222,u9temp_fifomodule222,u10carry_fifomodule222,u11carry_fifomodule222,empty_vc_buffer222_not_fifomodule2,u13temp_fifomodule222,u14temp_fifomodule222,u15carry_fifomodule222,u16carry_fifomodule222,u17res_fifomodule222,u18res_fifomodule222,write_ptr_ff_fifomodule222_0_not22,write_ptr_ff_fifomodule222_1_not22,b0wire_fifomodule222,b1wire_fifomodule222,u23temp_fifomodule222_not_fifomodule2,u23temp_fifomodule222,boutb_fifomodule222,bouta_fifomodule222,boutmain_fifomodule222,arst_value_fifomodule222;
	wire [33:0] flit22,flit221,flit222;
	wire [15:0] fifo_ff_fifomodule22,fifo_ff_fifomodule221,fifo_ff_fifomodule222;
	wire [1:0] write_ptr_ff_fifomodule22,read_ptr_ff_fifomodule22,next_write_ptr_fifomodule22,next_read_ptr_fifomodule22,fifo_ocup_fifomodule22,write_ptr_ff_fifomodule221,read_ptr_ff_fifomodule221,next_write_ptr_fifomodule221,next_read_ptr_fifomodule221,fifo_ocup_fifomodule221,write_ptr_ff_fifomodule222,read_ptr_ff_fifomodule222,next_write_ptr_fifomodule222,next_read_ptr_fifomodule222,fifo_ocup_fifomodule222;

	wire [110:0] from_input_req_in_jump_input_datapath3put_datapath3;
	wire [2:0] from_input_resp_input_datapath3;
	wire [110:0] to_output_req_in_jump_input_datapath3put_datapath3;
	wire [2:0] to_output_resp_input_datapath3;
	wire [1:0] vc_ch_act_in_input_datapath3;
	wire [1:0] vc_ch_act_out_input_datapath3;
	wire [2:0] i_input_datapath3;
	wire [2:0] j_input_datapath3;
	wire [0:1] _sv2v_jump_input_datapath3;

	wire req_in_jump_input_datapath3,req_out_jump_input_datapath3,xnor1resu_input_datapath3,xnor2resu_input_datapath3,and1resu_input_datapath3,cond1line_input_datapath3,req_in_jump_input_datapath3_not,and2resu_input_datapath3,xor1resu_input_datapath3,nand1resu_input_datapath33,xnor23resu_input_datapath3,and4resu_input_datapath3,write_flit3_vc_buffer3,norres_vc_buffer3_vc_buffer3,full_vc_buffer3,empty_vc_buffer3,error_vc_buffer3,read_flit3_vc_buffer3,locked_by_route_ff_vc_buffer3,next_locked_vc_buffer3,orres_vc_buffer3,or1res_vc_buffer3,or2res_vc_buffer3,finres1_vc_buffer3,andres1_vc_buffer3,full_vc_buffer3_not,locked_by_route_ff_vc_buffer3_not,thirdand_vc_buffer3,u1temp_fifomodule3,u2temp_fifomodule3,u4temp_fifomodule3,full_vc_buffer3_not_fifomodule,u7temp_fifomodule3,u9temp_fifomodule3,u10carry_fifomodule3,u11carry_fifomodule3,empty_vc_buffer3_not_fifomodule,u13temp_fifomodule3,u14temp_fifomodule3,u15carry_fifomodule3,u16carry_fifomodule3,u17res_fifomodule3,u18res_fifomodule3,write_ptr_ff_fifomodule3_0_not3,write_ptr_ff_fifomodule3_1_not3,b0wire_fifomodule3,b1wire_fifomodule3,u23temp_fifomodule3_not_fifomodule3,u23temp_fifomodule3,boutb_fifomodule3,bouta_fifomodule3,boutmain_fifomodule3,arst_value_fifomodule3,write_flit31_vc_buffer13,norres_vc_buffer31_vc_buffer1,full_vc_buffer31,empty_vc_buffer31,error_vc_buffer31,read_flit31_vc_buffer13,locked_by_route_ff_vc_buffer31,next_locked_vc_buffer31,orres_vc_buffer31,or1res_vc_buffer31,or2res_vc_buffer31,finres1_vc_buffer31,andres1_vc_buffer31,full_vc_buffer31_not1,locked_by_route_ff_vc_buffer31_not1,thirdand_vc_buffer31,u1temp_fifomodule31,u2temp_fifomodule31,u4temp_fifomodule31,full_vc_buffer31_not1_fifomodule1,u7temp_fifomodule31,u9temp_fifomodule31,u10carry_fifomodule31,u11carry_fifomodule31,empty_vc_buffer31_not_fifomodule1,u13temp_fifomodule31,u14temp_fifomodule31,u15carry_fifomodule31,u16carry_fifomodule31,u17res_fifomodule31,u18res_fifomodule31,write_ptr_ff_fifomodule31_0_not13,write_ptr_ff_fifomodule31_1_not13,b0wire_fifomodule31,b1wire_fifomodule31,u23temp_fifomodule31_not_fifomodule1,u23temp_fifomodule31,boutb_fifomodule31,bouta_fifomodule31,boutmain_fifomodule31,arst_value_fifomodule31,write_flit32_vc_buffer23,norres_vc_buffer32_vc_buffer2,full_vc_buffer32,empty_vc_buffer32,error_vc_buffer32,read_flit32_vc_buffer23,locked_by_route_ff_vc_buffer32,next_locked_vc_buffer32,orres_vc_buffer32,or1res_vc_buffer32,or2res_vc_buffer32,finres1_vc_buffer32,andres1_vc_buffer32,full_vc_buffer32_not2,locked_by_route_ff_vc_buffer32_not2,thirdand_vc_buffer32,u1temp_fifomodule32,u2temp_fifomodule32,u4temp_fifomodule32,full_vc_buffer32_not2_fifomodule2,u7temp_fifomodule32,u9temp_fifomodule32,u10carry_fifomodule32,u11carry_fifomodule32,empty_vc_buffer32_not_fifomodule2,u13temp_fifomodule32,u14temp_fifomodule32,u15carry_fifomodule32,u16carry_fifomodule32,u17res_fifomodule32,u18res_fifomodule32,write_ptr_ff_fifomodule32_0_not23,write_ptr_ff_fifomodule32_1_not23,b0wire_fifomodule32,b1wire_fifomodule32,u23temp_fifomodule32_not_fifomodule2,u23temp_fifomodule32,boutb_fifomodule32,bouta_fifomodule32,boutmain_fifomodule32,arst_value_fifomodule32;
	wire [33:0] flit3,flit31,flit32;
	wire [15:0] fifo_ff_fifomodule3,fifo_ff_fifomodule31,fifo_ff_fifomodule32;
	wire [1:0] write_ptr_ff_fifomodule3,read_ptr_ff_fifomodule3,next_write_ptr_fifomodule3,next_read_ptr_fifomodule3,fifo_ocup_fifomodule3,write_ptr_ff_fifomodule31,read_ptr_ff_fifomodule31,next_write_ptr_fifomodule31,next_read_ptr_fifomodule31,fifo_ocup_fifomodule31,write_ptr_ff_fifomodule32,read_ptr_ff_fifomodule32,next_write_ptr_fifomodule32,next_read_ptr_fifomodule32,fifo_ocup_fifomodule32;


	wire [110:0] from_input_req_in_jump_input_datapath4put_datapath4;
	wire [2:0] from_input_resp_input_datapath4;
	wire [110:0] to_output_req_in_jump_input_datapath4put_datapath4;
	wire [2:0] to_output_resp_input_datapath4;
	wire [1:0] vc_ch_act_in_input_datapath4;
	wire [1:0] vc_ch_act_out_input_datapath4;
	wire [2:0] i_input_datapath4;
	wire [2:0] j_input_datapath4;
	wire [0:1] _sv2v_jump_input_datapath4;

	wire req_in_jump_input_datapath4,req_out_jump_input_datapath4,xnor1resu_input_datapath4,xnor2resu_input_datapath4,and1resu_input_datapath4,cond1line_input_datapath4,req_in_jump_input_datapath4_not,and2resu_input_datapath4,xor1resu_input_datapath4,nand1resu_input_datapath44,xnor23resu_input_datapath4,and4resu_input_datapath4,write_flit4_vc_buffer4,norres_vc_buffer4_vc_buffer4,full_vc_buffer4,empty_vc_buffer4,error_vc_buffer4,read_flit4_vc_buffer4,locked_by_route_ff_vc_buffer4,next_locked_vc_buffer4,orres_vc_buffer4,or1res_vc_buffer4,or2res_vc_buffer4,finres1_vc_buffer4,andres1_vc_buffer4,full_vc_buffer4_not,locked_by_route_ff_vc_buffer4_not,thirdand_vc_buffer4,u1temp_fifomodule4,u2temp_fifomodule4,u4temp_fifomodule4,full_vc_buffer4_not_fifomodule,u7temp_fifomodule4,u9temp_fifomodule4,u10carry_fifomodule4,u11carry_fifomodule4,empty_vc_buffer4_not_fifomodule,u13temp_fifomodule4,u14temp_fifomodule4,u15carry_fifomodule4,u16carry_fifomodule4,u17res_fifomodule4,u18res_fifomodule4,write_ptr_ff_fifomodule4_0_not4,write_ptr_ff_fifomodule4_1_not4,b0wire_fifomodule4,b1wire_fifomodule4,u23temp_fifomodule4_not_fifomodule4,u23temp_fifomodule4,boutb_fifomodule4,bouta_fifomodule4,boutmain_fifomodule4,arst_value_fifomodule4,write_flit41_vc_buffer14,norres_vc_buffer41_vc_buffer1,full_vc_buffer41,empty_vc_buffer41,error_vc_buffer41,read_flit41_vc_buffer14,locked_by_route_ff_vc_buffer41,next_locked_vc_buffer41,orres_vc_buffer41,or1res_vc_buffer41,or2res_vc_buffer41,finres1_vc_buffer41,andres1_vc_buffer41,full_vc_buffer41_not1,locked_by_route_ff_vc_buffer41_not1,thirdand_vc_buffer41,u1temp_fifomodule41,u2temp_fifomodule41,u4temp_fifomodule41,full_vc_buffer41_not1_fifomodule1,u7temp_fifomodule41,u9temp_fifomodule41,u10carry_fifomodule41,u11carry_fifomodule41,empty_vc_buffer41_not_fifomodule1,u13temp_fifomodule41,u14temp_fifomodule41,u15carry_fifomodule41,u16carry_fifomodule41,u17res_fifomodule41,u18res_fifomodule41,write_ptr_ff_fifomodule41_0_not14,write_ptr_ff_fifomodule41_1_not14,b0wire_fifomodule41,b1wire_fifomodule41,u23temp_fifomodule41_not_fifomodule1,u23temp_fifomodule41,boutb_fifomodule41,bouta_fifomodule41,boutmain_fifomodule41,arst_value_fifomodule41,write_flit42_vc_buffer24,norres_vc_buffer42_vc_buffer2,full_vc_buffer42,empty_vc_buffer42,error_vc_buffer42,read_flit42_vc_buffer24,locked_by_route_ff_vc_buffer42,next_locked_vc_buffer42,orres_vc_buffer42,or1res_vc_buffer42,or2res_vc_buffer42,finres1_vc_buffer42,andres1_vc_buffer42,full_vc_buffer42_not2,locked_by_route_ff_vc_buffer42_not2,thirdand_vc_buffer42,u1temp_fifomodule42,u2temp_fifomodule42,u4temp_fifomodule42,full_vc_buffer42_not2_fifomodule2,u7temp_fifomodule42,u9temp_fifomodule42,u10carry_fifomodule42,u11carry_fifomodule42,empty_vc_buffer42_not_fifomodule2,u13temp_fifomodule42,u14temp_fifomodule42,u15carry_fifomodule42,u16carry_fifomodule42,u17res_fifomodule42,u18res_fifomodule42,write_ptr_ff_fifomodule42_0_not24,write_ptr_ff_fifomodule42_1_not24,b0wire_fifomodule42,b1wire_fifomodule42,u23temp_fifomodule42_not_fifomodule2,u23temp_fifomodule42,boutb_fifomodule42,bouta_fifomodule42,boutmain_fifomodule42,arst_value_fifomodule42;
	wire [33:0] flit4,flit41,flit42;
	wire [15:0] fifo_ff_fifomodule4,fifo_ff_fifomodule41,fifo_ff_fifomodule42;
	wire [1:0] write_ptr_ff_fifomodule4,read_ptr_ff_fifomodule4,next_write_ptr_fifomodule4,next_read_ptr_fifomodule4,fifo_ocup_fifomodule4,write_ptr_ff_fifomodule41,read_ptr_ff_fifomodule41,next_write_ptr_fifomodule41,next_read_ptr_fifomodule41,fifo_ocup_fifomodule41,write_ptr_ff_fifomodule42,read_ptr_ff_fifomodule42,next_write_ptr_fifomodule42,next_read_ptr_fifomodule42,fifo_ocup_fifomodule42;



//input router
    BUFX1 U0 ( .A(1'b0), .Y(next_rt_input_router[0]) );
    BUFX1 U1 ( .A(1'b0), .Y(next_rt_input_router[1]) );
    BUFX1 U2 ( .A(1'b0), .Y(next_rt_input_router[2]) );
    BUFX1 U3(.A(flit_input_router_req_i[3]), .Y(flit_input_router[3]));
	BUFX1 U4(.A(flit_input_router_req_i[4]), .Y(flit_input_router[4]));
	BUFX1 U5(.A(flit_input_router_req_i[5]), .Y(flit_input_router[5]));
	BUFX1 U6(.A(flit_input_router_req_i[6]), .Y(flit_input_router[6]));
	BUFX1 U7(.A(flit_input_router_req_i[7]), .Y(flit_input_router[7]));
	BUFX1 U8(.A(flit_input_router_req_i[8]), .Y(flit_input_router[8]));
	BUFX1 U9(.A(flit_input_router_req_i[9]), .Y(flit_input_router[9]));
	BUFX1 U10(.A(flit_input_router_req_i[10]), .Y(flit_input_router[10]));
	BUFX1 U11(.A(flit_input_router_req_i[11]), .Y(flit_input_router[11]));
	BUFX1 U12(.A(flit_input_router_req_i[12]), .Y(flit_input_router[12]));
	BUFX1 U13(.A(flit_input_router_req_i[13]), .Y(flit_input_router[13]));
	BUFX1 U14(.A(flit_input_router_req_i[14]), .Y(flit_input_router[14]));
	BUFX1 U15(.A(flit_input_router_req_i[15]), .Y(flit_input_router[15]));
	BUFX1 U16(.A(flit_input_router_req_i[16]), .Y(flit_input_router[16]));
	BUFX1 U17(.A(flit_input_router_req_i[17]), .Y(flit_input_router[17]));
	BUFX1 U18(.A(flit_input_router_req_i[18]), .Y(flit_input_router[18]));
	BUFX1 U19(.A(flit_input_router_req_i[19]), .Y(flit_input_router[19]));
	BUFX1 U20(.A(flit_input_router_req_i[20]), .Y(flit_input_router[20]));
	BUFX1 U21(.A(flit_input_router_req_i[21]), .Y(flit_input_router[21]));
	BUFX1 U22(.A(flit_input_router_req_i[22]), .Y(flit_input_router[22]));
	BUFX1 U23(.A(flit_input_router_req_i[23]), .Y(flit_input_router[23]));
	BUFX1 U24(.A(flit_input_router_req_i[24]), .Y(flit_input_router[24]));
	BUFX1 U25(.A(flit_input_router_req_i[25]), .Y(flit_input_router[25]));
	BUFX1 U26(.A(flit_input_router_req_i[26]), .Y(flit_input_router[26]));
	BUFX1 U27(.A(flit_input_router_req_i[27]), .Y(flit_input_router[27]));
	BUFX1 U28(.A(flit_input_router_req_i[28]), .Y(flit_input_router[28]));
	BUFX1 U29(.A(flit_input_router_req_i[29]), .Y(flit_input_router[29]));
	BUFX1 U30(.A(flit_input_router_req_i[30]), .Y(flit_input_router[30]));
	BUFX1 U31(.A(flit_input_router_req_i[31]), .Y(flit_input_router[31]));
	BUFX1 U32(.A(flit_input_router_req_i[32]), .Y(flit_input_router[32]));
	BUFX1 U33(.A(flit_input_router_req_i[33]), .Y(flit_input_router[33]));
	BUFX1 U34(.A(flit_input_router_req_i[34]), .Y(flit_input_router[34]));
	BUFX1 U35(.A(flit_input_router_req_i[35]), .Y(flit_input_router[35]));
	BUFX1 U36(.A(flit_input_router_req_i[36]), .Y(flit_input_router[36]));

    NOR2X1 U37 ( .IN1(flit_input_router[33]), .IN2(flit_input_router[32]), .QN(norres_1_input_router) );
    AND2X1 U38 ( .IN1(flit_input_router_req_i[0]), .IN2(norres_1_input_router), .Q(new_rt_input_router) );

    NOR2X1 U39 ( .IN1(flit_input_router[31]), .IN2(1'b0), .QN(norres_2_input_router) );
    NOR2X1 U40 ( .IN1(flit_input_router[30]), .IN2(1'b0), .QN(norres_3_input_router) );
    AND3X1 U41 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(norres_3_input_router), .Q(andfinres_input_router) );
    MUX21X1 U42 (.IN1(next_rt_input_router[0]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U43 (.IN1(next_rt_input_router[1]), .IN2(1'b0), .S(andfinres_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U44 (.IN1(next_rt_input_router[2]), .IN2(1'b1), .S(andfinres_input_router), .Q(next_rt_input_router[2]);
    INVX1 U45 ( .A(andfinres_input_router), .Y(invres1_input_router) );


    AND3X1 U46 ( .IN1(new_rt_input_router), .IN2(norres_2_input_router), .IN3(invres1_input_router), .Q(and2result_input_router) );
    MUX21X1 U47 (.IN1(next_rt_input_router[0]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U48 (.IN1(next_rt_input_router[1]), .IN2(1'b1), .S(and2result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U49 (.IN1(next_rt_input_router[2]), .IN2(1'b0), .S(and2result_input_router), .Q(next_rt_input_router[2]);
    INVX1 U50 ( .A(and2result_input_router), .Y(invres2_input_router) );

    AND3X1 U51 ( .IN1(new_rt_input_router), .IN2(invres1_input_router), .IN3(invres2_input_router), .Q(and3result_input_router) );
    AND2X1 U52 ( .IN1(flit_input_router[31]), .IN2(1'b1), .Q(and4result_input_router) );
    AND2X1 U53 ( .IN1(and4result_input_router), .IN2(and3result_input_router), .Q(and5result_input_router) );

    MUX21X1 U54 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router), .Q(next_rt_input_router[0]);
    MUX21X1 U55 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[1]);
    MUX21X1 U56 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router), .Q(next_rt_input_router[2]);

   	BUFX1 U57(.A(1'sb0), .Y(int_route_v[4:0][0]));
   	BUFX1 U58(.A(1'sb0), .Y(int_route_v[4:0][1]));
   	BUFX1 U59(.A(1'sb0), .Y(int_route_v[4:0][2]));
   	BUFX1 U60(.A(1'sb0), .Y(int_route_v[4:0][3]));
   	BUFX1 U61(.A(1'sb0), .Y(int_route_v[4:0][4]));

    NOR3X1 U62 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(norres_5_input_router) );
    AND2X1 U63 ( .IN1(norres_5_input_router), .IN2(new_rt_input_router), .Q(and6result_input_router) );
    MUX21X1 U64 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and6result_input_router), .Q(int_route_v[4:0][4]);

    NOR2X1 U65 ( .IN1(next_rt_input_router[1]), .IN2(next_rt_input_router[2]), .QN(and7result_input_router) );
    AND2X1 U66 ( .IN1(and7result_input_router), .IN2(next_rt_input_router[0]), .Y(orres1_input_router) );
    AND2X1 U67 ( .IN1(new_rt_input_router), .IN2(orres1_input_router), .Q(finand1_input_router) );
    MUX21X1 U68 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router), .Q(int_route_v[4:0][3]);

    NOR2X1 U69 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[2]), .Q(and8result_input_router) );
    AND2X1 U70 ( .IN1(and8result_input_router), .IN2(next_rt_input_router[1]), .Y(orres2_input_router) );
    AND2X1 U71 ( .IN1(new_rt_input_router), .IN2(orres2_input_router), .Q(finand2_input_router) );
    MUX21X1 U72 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router), .Q(int_route_v[4:0][2]);

    NOR2X1 U73 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and9result_input_router) );
    AND2X1 U74 ( .IN1(and9result_input_router), .IN2(next_rt_input_router[2]), .Y(orres3_input_router) );
    AND2X1 U75 ( .IN1(new_rt_input_router), .IN2(orres3_input_router), .Q(finand3_input_router) );
    MUX21X1 U76 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router), .Q(int_route_v[4:0][0]);

    AND2X1 U77 ( .IN1(next_rt_input_router[0]), .IN2(next_rt_input_router[1]), .Q(and10result_input_router) );
    INVX1 U78 ( .A(next_rt_input_router[2]), .Y(nextrt2not_input_router) );
    AND2X1 U79 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router), .Q(and11result_input_router) );
    MUX21X1 U80 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    INVX1 U81 ( .A(new_rt_input_router), .Y(new_rt_input_routernot) );
    AND2X1 U82 ( .IN1(new_rt_input_routernot), .IN2(flit_input_router_req_i[0]), .Q(secondAndc_input_router) );

    NOR3X1 U83 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(norres_5_input_router_2) );
    AND2X1 U84 ( .IN1(norres_5_input_router_2), .IN2(newsecondAndc_input_router_rt), .Q(and62result_input_router) );
    MUX21X1 U85 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(and62result_input_router), .Q(int_route_v[4:0][4]);

    NOR2X1 U86 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .QN(and7result_input_router2) );
    AND2X1 U87 ( .IN1(and7result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .Y(orres1_input_router2) );
    AND2X1 U88 ( .IN1(new_rt_input_routernot), .IN2(orres1_input_router2), .Q(finand1_input_router2) );
    MUX21X1 U89 (.IN1(int_route_v[4:0][3]), .IN2(1'sb1), .S(finand1_input_router2), .Q(int_route_v[4:0][3]);

    NOR2X1 U90 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Q(and8result_input_router2) );
    AND2X1 U91 ( .IN1(and8result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Y(orres2_input_router2) );
    AND2X1 U92 ( .IN1(new_rt_input_routernot), .IN2(orres2_input_router), .Q(finand2_input_router2) );
    MUX21X1 U93 (.IN1(int_route_v[4:0][2]), .IN2(1'sb1), .S(finand2_input_router2), .Q(int_route_v[4:0][2]);

    NOR2X1 U94 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and9result_input_router2) );
    AND2X1 U95 ( .IN1(and9result_input_router2), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(orres3_input_router2) );
    AND2X1 U96 ( .IN1(new_rt_input_routernot), .IN2(orres3_input_router2), .Q(finand3_input_router2) );
    MUX21X1 U97 (.IN1(int_route_v[4:0][0]), .IN2(1'sb1), .S(finand3_input_router2), .Q(int_route_v[4:0][0]);

    AND2X1 U98 ( .IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .Q(and10result_input_router2) );
    INVX1 U99 ( .A(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .Y(nextrt2not_input_router) );
    AND3X1 U100 ( .IN1(nextrt2not_input_router), .IN2(and10result_input_router2), .IN3(new_rt_input_routernot), .Q(and11result_input_router2) );
    MUX21X1 U101 (.IN1(int_route_v[4:0][1]), .IN2(1'sb1), .S(and11result_input_router), .Q(int_route_v[4:0][1]);

    DFFX2 U102 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U103 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U104 (.IN1(routing_table_ff_input_router[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[0]);
    MUX21X1 U105 (.IN1(routing_table_ff_input_router[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[1]);
    MUX21X1 U106 (.IN1(routing_table_ff_input_router[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[2]);
    MUX21X1 U107 (.IN1(routing_table_ff_input_router[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[3]);
    MUX21X1 U108 (.IN1(routing_table_ff_input_router[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[4]);
    MUX21X1 U109 (.IN1(routing_table_ff_input_router[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[5]);
    MUX21X1 U110 (.IN1(routing_table_ff_input_router[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[6]);
    MUX21X1 U111 (.IN1(routing_table_ff_input_router[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[7]);
    MUX21X1 U112 (.IN1(routing_table_ff_input_router[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router[8]);
    INVX1 U113 ( .A(arst_value), .Y(arst_valuenot_input_router) );
    AND2X1 U114 ( .IN1(new_rt_input_router), .IN2(arst_valuenot_input_router), .Q(finand3_input_router22) );
    MUX21X1 U115 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3]), .IN2(next_rt_input_router[0]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3]);
    MUX21X1 U116 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]), .IN2(next_rt_input_router[1]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+1]);
    MUX21X1 U117 (.IN1(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]), .IN2(next_rt_input_router[2]), .S(finand3_input_router22), .Q(routing_table_ff_input_router[flit_input_router_req_i[2]*3+2]);    

    BUFX1 U118 ( .A(1'b0), .Y(next_rt_input_router1[0]) );
    BUFX1 U119 ( .A(1'b0), .Y(next_rt_input_router1[1]) );
    BUFX1 U120 ( .A(1'b0), .Y(next_rt_input_router1[2]) );
    BUFX1 U121(.A(flit_input_router1_req_i[3]), .Y(flit_input_router1[3]));
    BUFX1 U122(.A(flit_input_router1_req_i[4]), .Y(flit_input_router1[4]));
    BUFX1 U123(.A(flit_input_router1_req_i[5]), .Y(flit_input_router1[5]));
    BUFX1 U124(.A(flit_input_router1_req_i[6]), .Y(flit_input_router1[6]));
    BUFX1 U125(.A(flit_input_router1_req_i[7]), .Y(flit_input_router1[7]));
    BUFX1 U126(.A(flit_input_router1_req_i[8]), .Y(flit_input_router1[8]));
    BUFX1 U127(.A(flit_input_router1_req_i[9]), .Y(flit_input_router1[9]));
    BUFX1 U128(.A(flit_input_router1_req_i[10]), .Y(flit_input_router1[10]));
    BUFX1 U129(.A(flit_input_router1_req_i[11]), .Y(flit_input_router1[11]));
    BUFX1 U130(.A(flit_input_router1_req_i[12]), .Y(flit_input_router1[12]));
    BUFX1 U131(.A(flit_input_router1_req_i[13]), .Y(flit_input_router1[13]));
    BUFX1 U132(.A(flit_input_router1_req_i[14]), .Y(flit_input_router1[14]));
    BUFX1 U133(.A(flit_input_router1_req_i[15]), .Y(flit_input_router1[15]));
    BUFX1 U134(.A(flit_input_router1_req_i[16]), .Y(flit_input_router1[16]));
    BUFX1 U135(.A(flit_input_router1_req_i[17]), .Y(flit_input_router1[17]));
    BUFX1 U136(.A(flit_input_router1_req_i[18]), .Y(flit_input_router1[18]));
    BUFX1 U137(.A(flit_input_router1_req_i[19]), .Y(flit_input_router1[19]));
    BUFX1 U138(.A(flit_input_router1_req_i[20]), .Y(flit_input_router1[20]));
    BUFX1 U139(.A(flit_input_router1_req_i[21]), .Y(flit_input_router1[21]));
    BUFX1 U140(.A(flit_input_router1_req_i[22]), .Y(flit_input_router1[22]));
    BUFX1 U141(.A(flit_input_router1_req_i[23]), .Y(flit_input_router1[23]));
    BUFX1 U142(.A(flit_input_router1_req_i[24]), .Y(flit_input_router1[24]));
    BUFX1 U143(.A(flit_input_router1_req_i[25]), .Y(flit_input_router1[25]));
    BUFX1 U144(.A(flit_input_router1_req_i[26]), .Y(flit_input_router1[26]));
    BUFX1 U145(.A(flit_input_router1_req_i[27]), .Y(flit_input_router1[27]));
    BUFX1 U146(.A(flit_input_router1_req_i[28]), .Y(flit_input_router1[28]));
    BUFX1 U147(.A(flit_input_router1_req_i[29]), .Y(flit_input_router1[29]));
    BUFX1 U148(.A(flit_input_router1_req_i[30]), .Y(flit_input_router1[30]));
    BUFX1 U149(.A(flit_input_router1_req_i[31]), .Y(flit_input_router1[31]));
    BUFX1 U150(.A(flit_input_router1_req_i[32]), .Y(flit_input_router1[32]));
    BUFX1 U151(.A(flit_input_router1_req_i[33]), .Y(flit_input_router1[33]));
    BUFX1 U152(.A(flit_input_router1_req_i[34]), .Y(flit_input_router1[34]));
    BUFX1 U153(.A(flit_input_router1_req_i[35]), .Y(flit_input_router1[35]));
    BUFX1 U154(.A(flit_input_router1_req_i[36]), .Y(flit_input_router1[36]));

    NOR2X1 U155 ( .IN1(flit_input_router1[33]), .IN2(flit_input_router1[32]), .QN(norres_1_input_router1) );
    AND2X1 U156 ( .IN1(flit_input_router1_req_i[0]), .IN2(norres_1_input_router1), .Q(new_rt_input_router1) );

    NOR2X1 U157 ( .IN1(flit_input_router1[31]), .IN2(1'b0), .QN(norres_2_input_router1) );
    NOR2X1 U158 ( .IN1(flit_input_router1[30]), .IN2(1'b0), .QN(norres_3_input_router1) );
    AND3X1 U159 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(norres_3_input_router1), .Q(andfinres_input_router1) );
    MUX21X1 U160 (.IN1(next_rt_input_router1[0]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U161 (.IN1(next_rt_input_router1[1]), .IN2(1'b0), .S(andfinres_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U162 (.IN1(next_rt_input_router1[2]), .IN2(1'b1), .S(andfinres_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U163 ( .A(andfinres_input_router1), .Y(invres1_input_router1) );


    AND3X1 U164 ( .IN1(new_rt_input_router1), .IN2(norres_2_input_router1), .IN3(invres1_input_router1), .Q(and2result_input_router1) );
    MUX21X1 U165 (.IN1(next_rt_input_router1[0]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U166 (.IN1(next_rt_input_router1[1]), .IN2(1'b1), .S(and2result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U167 (.IN1(next_rt_input_router1[2]), .IN2(1'b0), .S(and2result_input_router1), .Q(next_rt_input_router1[2]);
    INVX1 U168 ( .A(and2result_input_router1), .Y(invres2_input_router1) );

    AND3X1 U169 ( .IN1(new_rt_input_router1), .IN2(invres1_input_router1), .IN3(invres2_input_router1), .Q(and3result_input_router1) );
    AND2X1 U170 ( .IN1(flit_input_router1[31]), .IN2(1'b1), .Q(and4result_input_router1) );
    AND2X1 U171 ( .IN1(and4result_input_router1), .IN2(and3result_input_router1), .Q(and5result_input_router1) );

    MUX21X1 U172 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router1), .Q(next_rt_input_router1[0]);
    MUX21X1 U173 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[1]);
    MUX21X1 U174 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router1), .Q(next_rt_input_router1[2]);

    BUFX1 U175(.A(1'sb0), .Y(int_route_v[9:5][0]));
    BUFX1 U176(.A(1'sb0), .Y(int_route_v[9:5][1]));
    BUFX1 U177(.A(1'sb0), .Y(int_route_v[9:5][2]));
    BUFX1 U178(.A(1'sb0), .Y(int_route_v[9:5][3]));
    BUFX1 U179(.A(1'sb0), .Y(int_route_v[9:5][4]));

    NOR3X1 U180 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(norres_5_input_router1) );
    AND2X1 U181 ( .IN1(norres_5_input_router1), .IN2(new_rt_input_router1), .Q(and6result_input_router1) );
    MUX21X1 U182 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and6result_input_router1), .Q(int_route_v[9:5][4]);

    NOR2X1 U183 ( .IN1(next_rt_input_router1[1]), .IN2(next_rt_input_router1[2]), .QN(and7result_input_router1) );
    AND2X1 U184 ( .IN1(and7result_input_router1), .IN2(next_rt_input_router1[0]), .Y(orres1_input_router1) );
    AND2X1 U185 ( .IN1(new_rt_input_router1), .IN2(orres1_input_router1), .Q(finand1_input_router1) );
    MUX21X1 U186 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router1), .Q(int_route_v[9:5][3]);

    NOR2X1 U187 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[2]), .Q(and8result_input_router1) );
    AND2X1 U188 ( .IN1(and8result_input_router1), .IN2(next_rt_input_router1[1]), .Y(orres2_input_router1) );
    AND2X1 U189 ( .IN1(new_rt_input_router1), .IN2(orres2_input_router1), .Q(finand2_input_router1) );
    MUX21X1 U190 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router1), .Q(int_route_v[9:5][2]);

    NOR2X1 U191 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and9result_input_router1) );
    AND2X1 U192 ( .IN1(and9result_input_router1), .IN2(next_rt_input_router1[2]), .Y(orres3_input_router1) );
    AND2X1 U193 ( .IN1(new_rt_input_router1), .IN2(orres3_input_router1), .Q(finand3_input_router1) );
    MUX21X1 U194 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router1), .Q(int_route_v[9:5][0]);

    AND2X1 U195 ( .IN1(next_rt_input_router1[0]), .IN2(next_rt_input_router1[1]), .Q(and10result_input_router1) );
    INVX1 U196 ( .A(next_rt_input_router1[2]), .Y(nextrt2not_input_router11) );
    AND2X1 U197 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router1), .Q(and11result_input_router1) );
    MUX21X1 U198 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    INVX1 U199 ( .A(new_rt_input_router1), .Y(new_rt_input_router1not) );
    AND2X1 U200 ( .IN1(new_rt_input_router1not), .IN2(flit_input_router1_req_i[0]), .Q(secondAndc_input_router1) );

    NOR3X1 U201 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(norres_5_input_router1_2) );
    AND2X1 U202 ( .IN1(norres_5_input_router1_2), .IN2(newsecondAndc_input_router1_rt), .Q(and62result_input_router1) );
    MUX21X1 U203 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(and62result_input_router1), .Q(int_route_v[9:5][4]);

    NOR2X1 U204 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .QN(and7result_input_router12) );
    AND2X1 U205 ( .IN1(and7result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .Y(orres1_input_router12) );
    AND2X1 U206 ( .IN1(new_rt_input_router1not), .IN2(orres1_input_router12), .Q(finand1_input_router12) );
    MUX21X1 U207 (.IN1(int_route_v[9:5][3]), .IN2(1'sb1), .S(finand1_input_router12), .Q(int_route_v[9:5][3]);

    NOR2X1 U208 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Q(and8result_input_router12) );
    AND2X1 U209 ( .IN1(and8result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Y(orres2_input_router12) );
    AND2X1 U210 ( .IN1(new_rt_input_router1not), .IN2(orres2_input_router1), .Q(finand2_input_router12) );
    MUX21X1 U211 (.IN1(int_route_v[9:5][2]), .IN2(1'sb1), .S(finand2_input_router12), .Q(int_route_v[9:5][2]);

    NOR2X1 U212 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and9result_input_router12) );
    AND2X1 U213 ( .IN1(and9result_input_router12), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(orres3_input_router12) );
    AND2X1 U214 ( .IN1(new_rt_input_router1not), .IN2(orres3_input_router12), .Q(finand3_input_router12) );
    MUX21X1 U215 (.IN1(int_route_v[9:5][0]), .IN2(1'sb1), .S(finand3_input_router12), .Q(int_route_v[9:5][0]);

    AND2X1 U216 ( .IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .Q(and10result_input_router12) );
    INVX1 U217 ( .A(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .Y(nextrt2not_input_router11) );
    AND3X1 U218 ( .IN1(nextrt2not_input_router11), .IN2(and10result_input_router12), .IN3(new_rt_input_router1not), .Q(and11result_input_router12) );
    MUX21X1 U219 (.IN1(int_route_v[9:5][1]), .IN2(1'sb1), .S(and11result_input_router1), .Q(int_route_v[9:5][1]);

    DFFX2 U220 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U221 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U222 (.IN1(routing_table_ff_input_router1[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[0]);
    MUX21X1 U223 (.IN1(routing_table_ff_input_router1[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[1]);
    MUX21X1 U224 (.IN1(routing_table_ff_input_router1[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[2]);
    MUX21X1 U225 (.IN1(routing_table_ff_input_router1[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[3]);
    MUX21X1 U226 (.IN1(routing_table_ff_input_router1[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[4]);
    MUX21X1 U227 (.IN1(routing_table_ff_input_router1[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[5]);
    MUX21X1 U228 (.IN1(routing_table_ff_input_router1[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[6]);
    MUX21X1 U229 (.IN1(routing_table_ff_input_router1[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[7]);
    MUX21X1 U230 (.IN1(routing_table_ff_input_router1[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router1[8]);
    INVX1 U231 ( .A(arst_value), .Y(arst_valuenot_input_router1) );
    AND2X1 U232 ( .IN1(new_rt_input_router1), .IN2(arst_valuenot_input_router1), .Q(finand3_input_router122) );
    MUX21X1 U233 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]), .IN2(next_rt_input_router1[0]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3]);
    MUX21X1 U234 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]), .IN2(next_rt_input_router1[1]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+1]);
    MUX21X1 U235 (.IN1(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]), .IN2(next_rt_input_router1[2]), .S(finand3_input_router122), .Q(routing_table_ff_input_router1[flit_input_router1_req_i[2]*3+2]);


	BUFX1 U236 ( .A(1'b0), .Y(next_rt_input_router2[0]) );
    BUFX1 U237 ( .A(1'b0), .Y(next_rt_input_router2[1]) );
    BUFX1 U238 ( .A(1'b0), .Y(next_rt_input_router2[2]) );
    BUFX1 U239(.A(flit_input_router2_req_i[3]), .Y(flit_input_router2[3]));
    BUFX1 U240(.A(flit_input_router2_req_i[4]), .Y(flit_input_router2[4]));
    BUFX1 U241(.A(flit_input_router2_req_i[5]), .Y(flit_input_router2[5]));
    BUFX1 U242(.A(flit_input_router2_req_i[6]), .Y(flit_input_router2[6]));
    BUFX1 U243(.A(flit_input_router2_req_i[7]), .Y(flit_input_router2[7]));
    BUFX1 U244(.A(flit_input_router2_req_i[8]), .Y(flit_input_router2[8]));
    BUFX1 U245(.A(flit_input_router2_req_i[9]), .Y(flit_input_router2[9]));
    BUFX1 U246(.A(flit_input_router2_req_i[10]), .Y(flit_input_router2[10]));
    BUFX1 U247(.A(flit_input_router2_req_i[11]), .Y(flit_input_router2[11]));
    BUFX1 U248(.A(flit_input_router2_req_i[12]), .Y(flit_input_router2[12]));
    BUFX1 U249(.A(flit_input_router2_req_i[13]), .Y(flit_input_router2[13]));
    BUFX1 U250(.A(flit_input_router2_req_i[14]), .Y(flit_input_router2[14]));
    BUFX1 U251(.A(flit_input_router2_req_i[15]), .Y(flit_input_router2[15]));
    BUFX1 U252(.A(flit_input_router2_req_i[16]), .Y(flit_input_router2[16]));
    BUFX1 U253(.A(flit_input_router2_req_i[17]), .Y(flit_input_router2[17]));
    BUFX1 U254(.A(flit_input_router2_req_i[18]), .Y(flit_input_router2[18]));
    BUFX1 U255(.A(flit_input_router2_req_i[19]), .Y(flit_input_router2[19]));
    BUFX1 U256(.A(flit_input_router2_req_i[20]), .Y(flit_input_router2[20]));
    BUFX1 U257(.A(flit_input_router2_req_i[21]), .Y(flit_input_router2[21]));
    BUFX1 U258(.A(flit_input_router2_req_i[22]), .Y(flit_input_router2[22]));
    BUFX1 U259(.A(flit_input_router2_req_i[23]), .Y(flit_input_router2[23]));
    BUFX1 U260(.A(flit_input_router2_req_i[24]), .Y(flit_input_router2[24]));
    BUFX1 U261(.A(flit_input_router2_req_i[25]), .Y(flit_input_router2[25]));
    BUFX1 U262(.A(flit_input_router2_req_i[26]), .Y(flit_input_router2[26]));
    BUFX1 U263(.A(flit_input_router2_req_i[27]), .Y(flit_input_router2[27]));
    BUFX1 U264(.A(flit_input_router2_req_i[28]), .Y(flit_input_router2[28]));
    BUFX1 U265(.A(flit_input_router2_req_i[29]), .Y(flit_input_router2[29]));
    BUFX1 U266(.A(flit_input_router2_req_i[30]), .Y(flit_input_router2[30]));
    BUFX1 U267(.A(flit_input_router2_req_i[31]), .Y(flit_input_router2[31]));
    BUFX1 U268(.A(flit_input_router2_req_i[32]), .Y(flit_input_router2[32]));
    BUFX1 U269(.A(flit_input_router2_req_i[33]), .Y(flit_input_router2[33]));
    BUFX1 U270(.A(flit_input_router2_req_i[34]), .Y(flit_input_router2[34]));
    BUFX1 U271(.A(flit_input_router2_req_i[35]), .Y(flit_input_router2[35]));
    BUFX1 U272(.A(flit_input_router2_req_i[36]), .Y(flit_input_router2[36]));

    NOR2X1 U273 ( .IN1(flit_input_router2[33]), .IN2(flit_input_router2[32]), .QN(norres_1_input_router2) );
    AND2X1 U274 ( .IN1(flit_input_router2_req_i[0]), .IN2(norres_1_input_router2), .Q(new_rt_input_router2) );

    NOR2X1 U275 ( .IN1(flit_input_router2[31]), .IN2(1'b0), .QN(norres_2_input_router2) );
    NOR2X1 U276 ( .IN1(flit_input_router2[30]), .IN2(1'b0), .QN(norres_3_input_router2) );
    AND3X1 U277 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(norres_3_input_router2), .Q(andfinres_input_router2) );
    MUX21X1 U278 (.IN1(next_rt_input_router2[0]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U279 (.IN1(next_rt_input_router2[1]), .IN2(1'b0), .S(andfinres_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U280 (.IN1(next_rt_input_router2[2]), .IN2(1'b1), .S(andfinres_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U281 ( .A(andfinres_input_router2), .Y(invres1_input_router2) );


    AND3X1 U282 ( .IN1(new_rt_input_router2), .IN2(norres_2_input_router2), .IN3(invres1_input_router2), .Q(and2result_input_router2) );
    MUX21X1 U283 (.IN1(next_rt_input_router2[0]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U284 (.IN1(next_rt_input_router2[1]), .IN2(1'b1), .S(and2result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U285 (.IN1(next_rt_input_router2[2]), .IN2(1'b0), .S(and2result_input_router2), .Q(next_rt_input_router2[2]);
    INVX1 U286 ( .A(and2result_input_router2), .Y(invres2_input_router2) );

    AND3X1 U287 ( .IN1(new_rt_input_router2), .IN2(invres1_input_router2), .IN3(invres2_input_router2), .Q(and3result_input_router2) );
    AND2X1 U288 ( .IN1(flit_input_router2[31]), .IN2(1'b1), .Q(and4result_input_router2) );
    AND2X1 U289 ( .IN1(and4result_input_router2), .IN2(and3result_input_router2), .Q(and5result_input_router2) );

    MUX21X1 U290 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router2), .Q(next_rt_input_router2[0]);
    MUX21X1 U291 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[1]);
    MUX21X1 U292 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router2), .Q(next_rt_input_router2[2]);

    BUFX1 U293(.A(1'sb0), .Y(int_route_v[14:10][0]));
    BUFX1 U294(.A(1'sb0), .Y(int_route_v[14:10][1]));
    BUFX1 U295(.A(1'sb0), .Y(int_route_v[14:10][2]));
    BUFX1 U296(.A(1'sb0), .Y(int_route_v[14:10][3]));
    BUFX1 U297(.A(1'sb0), .Y(int_route_v[14:10][4]));

    NOR3X1 U298 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(norres_5_input_router2) );
    AND2X1 U299 ( .IN1(norres_5_input_router2), .IN2(new_rt_input_router2), .Q(and6result_input_router2) );
    MUX21X1 U300 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and6result_input_router2), .Q(int_route_v[14:10][4]);

    NOR2X1 U301 ( .IN1(next_rt_input_router2[1]), .IN2(next_rt_input_router2[2]), .QN(and7result_input_router22) );
    AND2X1 U302 ( .IN1(and7result_input_router22), .IN2(next_rt_input_router2[0]), .Y(orres1_input_router22) );
    AND2X1 U303 ( .IN1(new_rt_input_router2), .IN2(orres1_input_router22), .Q(finand1_input_router22) );
    MUX21X1 U304 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router22), .Q(int_route_v[14:10][3]);

    NOR2X1 U305 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[2]), .Q(and8result_input_router22) );
    AND2X1 U306 ( .IN1(and8result_input_router22), .IN2(next_rt_input_router2[1]), .Y(orres2_input_router22) );
    AND2X1 U307 ( .IN1(new_rt_input_router2), .IN2(orres2_input_router22), .Q(finand2_input_router22) );
    MUX21X1 U308 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router22), .Q(int_route_v[14:10][2]);

    NOR2X1 U309 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and9result_input_router22) );
    AND2X1 U310 ( .IN1(and9result_input_router22), .IN2(next_rt_input_router2[2]), .Y(orres3_input_router22) );
    AND2X1 U311 ( .IN1(new_rt_input_router2), .IN2(orres3_input_router22), .Q(finand3_input_router222) );
    MUX21X1 U312 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router222), .Q(int_route_v[14:10][0]);

    AND2X1 U313 ( .IN1(next_rt_input_router2[0]), .IN2(next_rt_input_router2[1]), .Q(and10result_input_router22) );
    INVX1 U314 ( .A(next_rt_input_router2[2]), .Y(nextrt2not_input_router22) );
    AND2X1 U315 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router22), .Q(and11result_input_router22) );
    MUX21X1 U316 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    INVX1 U317 ( .A(new_rt_input_router2), .Y(new_rt_input_router2not) );
    AND2X1 U318 ( .IN1(new_rt_input_router2not), .IN2(flit_input_router2_req_i[0]), .Q(secondAndc_input_router2) );

    NOR3X1 U319 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(norres_5_input_router2_2) );
    AND2X1 U320 ( .IN1(norres_5_input_router2_2), .IN2(newsecondAndc_input_router2_rt), .Q(and62result_input_router2) );
    MUX21X1 U321 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(and62result_input_router2), .Q(int_route_v[14:10][4]);

    NOR2X1 U322 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .QN(and7result_input_router222) );
    AND2X1 U323 ( .IN1(and7result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .Y(orres1_input_router222) );
    AND2X1 U324 ( .IN1(new_rt_input_router2not), .IN2(orres1_input_router222), .Q(finand1_input_router222) );
    MUX21X1 U325 (.IN1(int_route_v[14:10][3]), .IN2(1'sb1), .S(finand1_input_router222), .Q(int_route_v[14:10][3]);

    NOR2X1 U326 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Q(and8result_input_router222) );
    AND2X1 U327 ( .IN1(and8result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Y(orres2_input_router222) );
    AND2X1 U328 ( .IN1(new_rt_input_router2not), .IN2(orres2_input_router22), .Q(finand2_input_router222) );
    MUX21X1 U329 (.IN1(int_route_v[14:10][2]), .IN2(1'sb1), .S(finand2_input_router222), .Q(int_route_v[14:10][2]);

    NOR2X1 U330 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and9result_input_router222) );
    AND2X1 U331 ( .IN1(and9result_input_router222), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(orres3_input_router222) );
    AND2X1 U332 ( .IN1(new_rt_input_router2not), .IN2(orres3_input_router222), .Q(finand3_input_router2222) );
    MUX21X1 U333 (.IN1(int_route_v[14:10][0]), .IN2(1'sb1), .S(finand3_input_router2222), .Q(int_route_v[14:10][0]);

    AND2X1 U334 ( .IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .Q(and10result_input_router222) );
    INVX1 U335 ( .A(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .Y(nextrt2not_input_router22) );
    AND3X1 U336 ( .IN1(nextrt2not_input_router22), .IN2(and10result_input_router222), .IN3(new_rt_input_router2not), .Q(and11result_input_router222) );
    MUX21X1 U337 (.IN1(int_route_v[14:10][1]), .IN2(1'sb1), .S(and11result_input_router22), .Q(int_route_v[14:10][1]);

    DFFX2 U338 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U339 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U340 (.IN1(routing_table_ff_input_router2[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[0]);
    MUX21X1 U341 (.IN1(routing_table_ff_input_router2[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[1]);
    MUX21X1 U342 (.IN1(routing_table_ff_input_router2[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[2]);
    MUX21X1 U343 (.IN1(routing_table_ff_input_router2[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[3]);
    MUX21X1 U344 (.IN1(routing_table_ff_input_router2[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[4]);
    MUX21X1 U345 (.IN1(routing_table_ff_input_router2[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[5]);
    MUX21X1 U346 (.IN1(routing_table_ff_input_router2[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[6]);
    MUX21X1 U347 (.IN1(routing_table_ff_input_router2[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[7]);
    MUX21X1 U348 (.IN1(routing_table_ff_input_router2[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router2[8]);
    INVX1 U349 ( .A(arst_value), .Y(arst_valuenot_input_router2) );
    AND2X1 U350 ( .IN1(new_rt_input_router2), .IN2(arst_valuenot_input_router2), .Q(finand3_input_router22222) );
    MUX21X1 U351 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]), .IN2(next_rt_input_router2[0]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3]);
    MUX21X1 U352 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]), .IN2(next_rt_input_router2[1]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+1]);
    MUX21X1 U353 (.IN1(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]), .IN2(next_rt_input_router2[2]), .S(finand3_input_router22222), .Q(routing_table_ff_input_router2[flit_input_router2_req_i[2]*3+2]); 

    BUFX1 U354 ( .A(1'b0), .Y(next_rt_input_router3[0]) );
    BUFX1 U355 ( .A(1'b0), .Y(next_rt_input_router3[1]) );
    BUFX1 U356 ( .A(1'b0), .Y(next_rt_input_router3[2]) );
    BUFX1 U357(.A(flit_input_router3_req_i[3]), .Y(flit_input_router3[3]));
    BUFX1 U358(.A(flit_input_router3_req_i[4]), .Y(flit_input_router3[4]));
    BUFX1 U359(.A(flit_input_router3_req_i[5]), .Y(flit_input_router3[5]));
    BUFX1 U360(.A(flit_input_router3_req_i[6]), .Y(flit_input_router3[6]));
    BUFX1 U361(.A(flit_input_router3_req_i[7]), .Y(flit_input_router3[7]));
    BUFX1 U362(.A(flit_input_router3_req_i[8]), .Y(flit_input_router3[8]));
    BUFX1 U363(.A(flit_input_router3_req_i[9]), .Y(flit_input_router3[9]));
    BUFX1 U364(.A(flit_input_router3_req_i[10]), .Y(flit_input_router3[10]));
    BUFX1 U365(.A(flit_input_router3_req_i[11]), .Y(flit_input_router3[11]));
    BUFX1 U366(.A(flit_input_router3_req_i[12]), .Y(flit_input_router3[12]));
    BUFX1 U367(.A(flit_input_router3_req_i[13]), .Y(flit_input_router3[13]));
    BUFX1 U368(.A(flit_input_router3_req_i[14]), .Y(flit_input_router3[14]));
    BUFX1 U369(.A(flit_input_router3_req_i[15]), .Y(flit_input_router3[15]));
    BUFX1 U370(.A(flit_input_router3_req_i[16]), .Y(flit_input_router3[16]));
    BUFX1 U371(.A(flit_input_router3_req_i[17]), .Y(flit_input_router3[17]));
    BUFX1 U372(.A(flit_input_router3_req_i[18]), .Y(flit_input_router3[18]));
    BUFX1 U373(.A(flit_input_router3_req_i[19]), .Y(flit_input_router3[19]));
    BUFX1 U374(.A(flit_input_router3_req_i[20]), .Y(flit_input_router3[20]));
    BUFX1 U375(.A(flit_input_router3_req_i[21]), .Y(flit_input_router3[21]));
    BUFX1 U376(.A(flit_input_router3_req_i[22]), .Y(flit_input_router3[22]));
    BUFX1 U377(.A(flit_input_router3_req_i[23]), .Y(flit_input_router3[23]));
    BUFX1 U378(.A(flit_input_router3_req_i[24]), .Y(flit_input_router3[24]));
    BUFX1 U379(.A(flit_input_router3_req_i[25]), .Y(flit_input_router3[25]));
    BUFX1 U380(.A(flit_input_router3_req_i[26]), .Y(flit_input_router3[26]));
    BUFX1 U381(.A(flit_input_router3_req_i[27]), .Y(flit_input_router3[27]));
    BUFX1 U382(.A(flit_input_router3_req_i[28]), .Y(flit_input_router3[28]));
    BUFX1 U383(.A(flit_input_router3_req_i[29]), .Y(flit_input_router3[29]));
    BUFX1 U384(.A(flit_input_router3_req_i[30]), .Y(flit_input_router3[30]));
    BUFX1 U385(.A(flit_input_router3_req_i[31]), .Y(flit_input_router3[31]));
    BUFX1 U386(.A(flit_input_router3_req_i[32]), .Y(flit_input_router3[32]));
    BUFX1 U387(.A(flit_input_router3_req_i[33]), .Y(flit_input_router3[33]));
    BUFX1 U388(.A(flit_input_router3_req_i[34]), .Y(flit_input_router3[34]));
    BUFX1 U389(.A(flit_input_router3_req_i[35]), .Y(flit_input_router3[35]));
    BUFX1 U390(.A(flit_input_router3_req_i[36]), .Y(flit_input_router3[36]));

    NOR2X1 U391 ( .IN1(flit_input_router3[33]), .IN2(flit_input_router3[32]), .QN(norres_1_input_router3) );
    AND2X1 U392 ( .IN1(flit_input_router3_req_i[0]), .IN2(norres_1_input_router3), .Q(new_rt_input_router3) );

    NOR2X1 U393 ( .IN1(flit_input_router3[31]), .IN2(1'b0), .QN(norres_2_input_router3) );
    NOR2X1 U394 ( .IN1(flit_input_router3[30]), .IN2(1'b0), .QN(norres_3_input_router3) );
    AND3X1 U395 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(norres_3_input_router3), .Q(andfinres_input_router3) );
    MUX21X1 U396 (.IN1(next_rt_input_router3[0]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U397 (.IN1(next_rt_input_router3[1]), .IN2(1'b0), .S(andfinres_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U398 (.IN1(next_rt_input_router3[2]), .IN2(1'b1), .S(andfinres_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U399 ( .A(andfinres_input_router3), .Y(invres1_input_router3) );


    AND3X1 U400 ( .IN1(new_rt_input_router3), .IN2(norres_2_input_router3), .IN3(invres1_input_router3), .Q(and2result_input_router3) );
    MUX21X1 U401 (.IN1(next_rt_input_router3[0]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U402 (.IN1(next_rt_input_router3[1]), .IN2(1'b1), .S(and2result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U403 (.IN1(next_rt_input_router3[2]), .IN2(1'b0), .S(and2result_input_router3), .Q(next_rt_input_router3[2]);
    INVX1 U404 ( .A(and2result_input_router3), .Y(invres2_input_router3) );

    AND3X1 U405 ( .IN1(new_rt_input_router3), .IN2(invres1_input_router3), .IN3(invres2_input_router3), .Q(and3result_input_router3) );
    AND2X1 U406 ( .IN1(flit_input_router3[31]), .IN2(1'b1), .Q(and4result_input_router3) );
    AND2X1 U407 ( .IN1(and4result_input_router3), .IN2(and3result_input_router3), .Q(and5result_input_router3) );

    MUX21X1 U408 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router3), .Q(next_rt_input_router3[0]);
    MUX21X1 U409 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[1]);
    MUX21X1 U410 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router3), .Q(next_rt_input_router3[2]);

    BUFX1 U411(.A(1'sb0), .Y(int_route_v[19:15][0]));
    BUFX1 U412(.A(1'sb0), .Y(int_route_v[19:15][1]));
    BUFX1 U413(.A(1'sb0), .Y(int_route_v[19:15][2]));
    BUFX1 U414(.A(1'sb0), .Y(int_route_v[19:15][3]));
    BUFX1 U415(.A(1'sb0), .Y(int_route_v[19:15][4]));

    NOR3X1 U416 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(norres_5_input_router3) );
    AND2X1 U417 ( .IN1(norres_5_input_router3), .IN2(new_rt_input_router3), .Q(and6result_input_router3) );
    MUX21X1 U418 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and6result_input_router3), .Q(int_route_v[19:15][4]);

    NOR2X1 U419 ( .IN1(next_rt_input_router3[1]), .IN2(next_rt_input_router3[2]), .QN(and7result_input_router3) );
    AND2X1 U420 ( .IN1(and7result_input_router3), .IN2(next_rt_input_router3[0]), .Y(orres1_input_router3) );
    AND2X1 U421 ( .IN1(new_rt_input_router3), .IN2(orres1_input_router3), .Q(finand1_input_router3) );
    MUX21X1 U422 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router3), .Q(int_route_v[19:15][3]);

    NOR2X1 U423 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[2]), .Q(and8result_input_router3) );
    AND2X1 U424 ( .IN1(and8result_input_router3), .IN2(next_rt_input_router3[1]), .Y(orres2_input_router3) );
    AND2X1 U425 ( .IN1(new_rt_input_router3), .IN2(orres2_input_router3), .Q(finand2_input_router3) );
    MUX21X1 U426 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router3), .Q(int_route_v[19:15][2]);

    NOR2X1 U427 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and9result_input_router3) );
    AND2X1 U428 ( .IN1(and9result_input_router3), .IN2(next_rt_input_router3[2]), .Y(orres3_input_router3) );
    AND2X1 U429 ( .IN1(new_rt_input_router3), .IN2(orres3_input_router3), .Q(finand3_input_router3) );
    MUX21X1 U430 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router3), .Q(int_route_v[19:15][0]);

    AND2X1 U431 ( .IN1(next_rt_input_router3[0]), .IN2(next_rt_input_router3[1]), .Q(and10result_input_router3) );
    INVX1 U432 ( .A(next_rt_input_router3[2]), .Y(nextrt2not_input_router33) );
    AND2X1 U433 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router3), .Q(and11result_input_router3) );
    MUX21X1 U434 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    INVX1 U435 ( .A(new_rt_input_router3), .Y(new_rt_input_router3not) );
    AND2X1 U436 ( .IN1(new_rt_input_router3not), .IN2(flit_input_router3_req_i[0]), .Q(secondAndc_input_router3) );

    NOR3X1 U437 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(norres_5_input_router3_2) );
    AND2X1 U438 ( .IN1(norres_5_input_router3_2), .IN2(newsecondAndc_input_router3_rt), .Q(and62result_input_router3) );
    MUX21X1 U439 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(and62result_input_router3), .Q(int_route_v[19:15][4]);

    NOR2X1 U440 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .QN(and7result_input_router32) );
    AND2X1 U441 ( .IN1(and7result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .Y(orres1_input_router32) );
    AND2X1 U442 ( .IN1(new_rt_input_router3not), .IN2(orres1_input_router32), .Q(finand1_input_router32) );
    MUX21X1 U443 (.IN1(int_route_v[19:15][3]), .IN2(1'sb1), .S(finand1_input_router32), .Q(int_route_v[19:15][3]);

    NOR2X1 U444 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Q(and8result_input_router32) );
    AND2X1 U445 ( .IN1(and8result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Y(orres2_input_router32) );
    AND2X1 U446 ( .IN1(new_rt_input_router3not), .IN2(orres2_input_router3), .Q(finand2_input_router32) );
    MUX21X1 U447 (.IN1(int_route_v[19:15][2]), .IN2(1'sb1), .S(finand2_input_router32), .Q(int_route_v[19:15][2]);

    NOR2X1 U448 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and9result_input_router32) );
    AND2X1 U449 ( .IN1(and9result_input_router32), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(orres3_input_router32) );
    AND2X1 U450 ( .IN1(new_rt_input_router3not), .IN2(orres3_input_router32), .Q(finand3_input_router32) );
    MUX21X1 U451 (.IN1(int_route_v[19:15][0]), .IN2(1'sb1), .S(finand3_input_router32), .Q(int_route_v[19:15][0]);

    AND2X1 U452 ( .IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .Q(and10result_input_router32) );
    INVX1 U453 ( .A(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .Y(nextrt2not_input_router33) );
    AND3X1 U454 ( .IN1(nextrt2not_input_router33), .IN2(and10result_input_router32), .IN3(new_rt_input_router3not), .Q(and11result_input_router32) );
    MUX21X1 U455 (.IN1(int_route_v[19:15][1]), .IN2(1'sb1), .S(and11result_input_router3), .Q(int_route_v[19:15][1]);

    DFFX2 U456 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U457 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U458 (.IN1(routing_table_ff_input_router3[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[0]);
    MUX21X1 U459 (.IN1(routing_table_ff_input_router3[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[1]);
    MUX21X1 U460 (.IN1(routing_table_ff_input_router3[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[2]);
    MUX21X1 U461 (.IN1(routing_table_ff_input_router3[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[3]);
    MUX21X1 U462 (.IN1(routing_table_ff_input_router3[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[4]);
    MUX21X1 U463 (.IN1(routing_table_ff_input_router3[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[5]);
    MUX21X1 U464 (.IN1(routing_table_ff_input_router3[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[6]);
    MUX21X1 U465 (.IN1(routing_table_ff_input_router3[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[7]);
    MUX21X1 U466 (.IN1(routing_table_ff_input_router3[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router3[8]);
    INVX1 U467 ( .A(arst_value), .Y(arst_valuenot_input_router3) );
    AND2X1 U468 ( .IN1(new_rt_input_router3), .IN2(arst_valuenot_input_router3), .Q(finand3_input_router322) );
    MUX21X1 U469 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]), .IN2(next_rt_input_router3[0]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3]);
    MUX21X1 U470 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]), .IN2(next_rt_input_router3[1]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+1]);
    MUX21X1 U471 (.IN1(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]), .IN2(next_rt_input_router3[2]), .S(finand3_input_router322), .Q(routing_table_ff_input_router3[flit_input_router3_req_i[2]*3+2]);

    BUFX1 U472 ( .A(1'b0), .Y(next_rt_input_router4[0]) );
    BUFX1 U473 ( .A(1'b0), .Y(next_rt_input_router4[1]) );
    BUFX1 U474 ( .A(1'b0), .Y(next_rt_input_router4[2]) );
    BUFX1 U475(.A(flit_input_router4_req_i[3]), .Y(flit_input_router4[3]));
    BUFX1 U476(.A(flit_input_router4_req_i[4]), .Y(flit_input_router4[4]));
    BUFX1 U477(.A(flit_input_router4_req_i[5]), .Y(flit_input_router4[5]));
    BUFX1 U478(.A(flit_input_router4_req_i[6]), .Y(flit_input_router4[6]));
    BUFX1 U479(.A(flit_input_router4_req_i[7]), .Y(flit_input_router4[7]));
    BUFX1 U480(.A(flit_input_router4_req_i[8]), .Y(flit_input_router4[8]));
    BUFX1 U481(.A(flit_input_router4_req_i[9]), .Y(flit_input_router4[9]));
    BUFX1 U482(.A(flit_input_router4_req_i[10]), .Y(flit_input_router4[10]));
    BUFX1 U483(.A(flit_input_router4_req_i[11]), .Y(flit_input_router4[11]));
    BUFX1 U484(.A(flit_input_router4_req_i[12]), .Y(flit_input_router4[12]));
    BUFX1 U485(.A(flit_input_router4_req_i[13]), .Y(flit_input_router4[13]));
    BUFX1 U486(.A(flit_input_router4_req_i[14]), .Y(flit_input_router4[14]));
    BUFX1 U487(.A(flit_input_router4_req_i[15]), .Y(flit_input_router4[15]));
    BUFX1 U488(.A(flit_input_router4_req_i[16]), .Y(flit_input_router4[16]));
    BUFX1 U489(.A(flit_input_router4_req_i[17]), .Y(flit_input_router4[17]));
    BUFX1 U490(.A(flit_input_router4_req_i[18]), .Y(flit_input_router4[18]));
    BUFX1 U491(.A(flit_input_router4_req_i[19]), .Y(flit_input_router4[19]));
    BUFX1 U492(.A(flit_input_router4_req_i[20]), .Y(flit_input_router4[20]));
    BUFX1 U493(.A(flit_input_router4_req_i[21]), .Y(flit_input_router4[21]));
    BUFX1 U494(.A(flit_input_router4_req_i[22]), .Y(flit_input_router4[22]));
    BUFX1 U495(.A(flit_input_router4_req_i[23]), .Y(flit_input_router4[23]));
    BUFX1 U496(.A(flit_input_router4_req_i[24]), .Y(flit_input_router4[24]));
    BUFX1 U497(.A(flit_input_router4_req_i[25]), .Y(flit_input_router4[25]));
    BUFX1 U498(.A(flit_input_router4_req_i[26]), .Y(flit_input_router4[26]));
    BUFX1 U499(.A(flit_input_router4_req_i[27]), .Y(flit_input_router4[27]));
    BUFX1 U500(.A(flit_input_router4_req_i[28]), .Y(flit_input_router4[28]));
    BUFX1 U501(.A(flit_input_router4_req_i[29]), .Y(flit_input_router4[29]));
    BUFX1 U502(.A(flit_input_router4_req_i[30]), .Y(flit_input_router4[30]));
    BUFX1 U503(.A(flit_input_router4_req_i[31]), .Y(flit_input_router4[31]));
    BUFX1 U504(.A(flit_input_router4_req_i[32]), .Y(flit_input_router4[32]));
    BUFX1 U505(.A(flit_input_router4_req_i[33]), .Y(flit_input_router4[33]));
    BUFX1 U506(.A(flit_input_router4_req_i[34]), .Y(flit_input_router4[34]));
    BUFX1 U507(.A(flit_input_router4_req_i[35]), .Y(flit_input_router4[35]));
    BUFX1 U508(.A(flit_input_router4_req_i[36]), .Y(flit_input_router4[36]));

    NOR2X1 U509 ( .IN1(flit_input_router4[33]), .IN2(flit_input_router4[32]), .QN(norres_1_input_router4) );
    AND2X1 U510 ( .IN1(flit_input_router4_req_i[0]), .IN2(norres_1_input_router4), .Q(new_rt_input_router4) );

    NOR2X1 U511 ( .IN1(flit_input_router4[31]), .IN2(1'b0), .QN(norres_2_input_router4) );
    NOR2X1 U512 ( .IN1(flit_input_router4[30]), .IN2(1'b0), .QN(norres_3_input_router4) );
    AND3X1 U513 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(norres_3_input_router4), .Q(andfinres_input_router4) );
    MUX21X1 U514 (.IN1(next_rt_input_router4[0]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U515 (.IN1(next_rt_input_router4[1]), .IN2(1'b0), .S(andfinres_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U516 (.IN1(next_rt_input_router4[2]), .IN2(1'b1), .S(andfinres_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U517 ( .A(andfinres_input_router4), .Y(invres1_input_router4) );


    AND3X1 U518 ( .IN1(new_rt_input_router4), .IN2(norres_2_input_router4), .IN3(invres1_input_router4), .Q(and2result_input_router4) );
    MUX21X1 U519 (.IN1(next_rt_input_router4[0]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U520 (.IN1(next_rt_input_router4[1]), .IN2(1'b1), .S(and2result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U521 (.IN1(next_rt_input_router4[2]), .IN2(1'b0), .S(and2result_input_router4), .Q(next_rt_input_router4[2]);
    INVX1 U522 ( .A(and2result_input_router4), .Y(invres2_input_router4) );

    AND3X1 U523 ( .IN1(new_rt_input_router4), .IN2(invres1_input_router4), .IN3(invres2_input_router4), .Q(and3result_input_router4) );
    AND2X1 U524 ( .IN1(flit_input_router4[31]), .IN2(1'b1), .Q(and4result_input_router4) );
    AND2X1 U525 ( .IN1(and4result_input_router4), .IN2(and3result_input_router4), .Q(and5result_input_router4) );

    MUX21X1 U526 (.IN1(1'b0), .IN2(1'b1), .S(and5result_input_router4), .Q(next_rt_input_router4[0]);
    MUX21X1 U527 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[1]);
    MUX21X1 U528 (.IN1(1'b0), .IN2(1'b0), .S(and5result_input_router4), .Q(next_rt_input_router4[2]);

    BUFX1 U529(.A(1'sb0), .Y(int_route_v[24:20][0]));
    BUFX1 U530(.A(1'sb0), .Y(int_route_v[24:20][1]));
    BUFX1 U531(.A(1'sb0), .Y(int_route_v[24:20][2]));
    BUFX1 U532(.A(1'sb0), .Y(int_route_v[24:20][3]));
    BUFX1 U533(.A(1'sb0), .Y(int_route_v[24:20][4]));

    NOR3X1 U534 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(norres_5_input_router4) );
    AND2X1 U535 ( .IN1(norres_5_input_router4), .IN2(new_rt_input_router4), .Q(and6result_input_router4) );
    MUX21X1 U536 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and6result_input_router4), .Q(int_route_v[24:20][4]);

    NOR2X1 U537 ( .IN1(next_rt_input_router4[1]), .IN2(next_rt_input_router4[2]), .QN(and7result_input_router4) );
    AND2X1 U538 ( .IN1(and7result_input_router4), .IN2(next_rt_input_router4[0]), .Y(orres1_input_router4) );
    AND2X1 U539 ( .IN1(new_rt_input_router4), .IN2(orres1_input_router4), .Q(finand1_input_router4) );
    MUX21X1 U540 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router4), .Q(int_route_v[24:20][3]);

    NOR2X1 U541 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[2]), .Q(and8result_input_router4) );
    AND2X1 U542 ( .IN1(and8result_input_router4), .IN2(next_rt_input_router4[1]), .Y(orres2_input_router4) );
    AND2X1 U543 ( .IN1(new_rt_input_router4), .IN2(orres2_input_router4), .Q(finand2_input_router4) );
    MUX21X1 U544 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router4), .Q(int_route_v[24:20][2]);

    NOR2X1 U545 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and9result_input_router4) );
    AND2X1 U546 ( .IN1(and9result_input_router4), .IN2(next_rt_input_router4[2]), .Y(orres3_input_router4) );
    AND2X1 U547 ( .IN1(new_rt_input_router4), .IN2(orres3_input_router4), .Q(finand3_input_router4) );
    MUX21X1 U548 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router4), .Q(int_route_v[24:20][0]);

    AND2X1 U549 ( .IN1(next_rt_input_router4[0]), .IN2(next_rt_input_router4[1]), .Q(and10result_input_router4) );
    INVX1 U550 ( .A(next_rt_input_router4[2]), .Y(nextrt2not_input_router44) );
    AND2X1 U551 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router4), .Q(and11result_input_router4) );
    MUX21X1 U552 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    INVX1 U553 ( .A(new_rt_input_router4), .Y(new_rt_input_router4not) );
    AND2X1 U554 ( .IN1(new_rt_input_router4not), .IN2(flit_input_router4_req_i[0]), .Q(secondAndc_input_router4) );

    NOR3X1 U555 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(norres_5_input_router4_2) );
    AND2X1 U556 ( .IN1(norres_5_input_router4_2), .IN2(newsecondAndc_input_router4_rt), .Q(and62result_input_router4) );
    MUX21X1 U557 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(and62result_input_router4), .Q(int_route_v[24:20][4]);

    NOR2X1 U558 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .QN(and7result_input_router42) );
    AND2X1 U559 ( .IN1(and7result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .Y(orres1_input_router42) );
    AND2X1 U560 ( .IN1(new_rt_input_router4not), .IN2(orres1_input_router42), .Q(finand1_input_router42) );
    MUX21X1 U561 (.IN1(int_route_v[24:20][3]), .IN2(1'sb1), .S(finand1_input_router42), .Q(int_route_v[24:20][3]);

    NOR2X1 U562 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Q(and8result_input_router42) );
    AND2X1 U563 ( .IN1(and8result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Y(orres2_input_router42) );
    AND2X1 U564 ( .IN1(new_rt_input_router4not), .IN2(orres2_input_router4), .Q(finand2_input_router42) );
    MUX21X1 U565 (.IN1(int_route_v[24:20][2]), .IN2(1'sb1), .S(finand2_input_router42), .Q(int_route_v[24:20][2]);

    NOR2X1 U566 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and9result_input_router42) );
    AND2X1 U567 ( .IN1(and9result_input_router42), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(orres3_input_router42) );
    AND2X1 U568 ( .IN1(new_rt_input_router4not), .IN2(orres3_input_router42), .Q(finand3_input_router42) );
    MUX21X1 U569 (.IN1(int_route_v[24:20][0]), .IN2(1'sb1), .S(finand3_input_router42), .Q(int_route_v[24:20][0]);

    AND2X1 U570 ( .IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .Q(and10result_input_router42) );
    INVX1 U571 ( .A(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .Y(nextrt2not_input_router44) );
    AND3X1 U572 ( .IN1(nextrt2not_input_router44), .IN2(and10result_input_router42), .IN3(new_rt_input_router4not), .Q(and11result_input_router42) );
    MUX21X1 U573 (.IN1(int_route_v[24:20][1]), .IN2(1'sb1), .S(and11result_input_router4), .Q(int_route_v[24:20][1]);

    DFFX2 U574 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U575 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U576 (.IN1(routing_table_ff_input_router4[0]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[0]);
    MUX21X1 U577 (.IN1(routing_table_ff_input_router4[1]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[1]);
    MUX21X1 U578 (.IN1(routing_table_ff_input_router4[2]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[2]);
    MUX21X1 U579 (.IN1(routing_table_ff_input_router4[3]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[3]);
    MUX21X1 U580 (.IN1(routing_table_ff_input_router4[4]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[4]);
    MUX21X1 U581 (.IN1(routing_table_ff_input_router4[5]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[5]);
    MUX21X1 U582 (.IN1(routing_table_ff_input_router4[6]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[6]);
    MUX21X1 U583 (.IN1(routing_table_ff_input_router4[7]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[7]);
    MUX21X1 U584 (.IN1(routing_table_ff_input_router4[8]), .IN2(1'sb0), .S(arst_value), .Q(routing_table_ff_input_router4[8]);
    INVX1 U585 ( .A(arst_value), .Y(arst_valuenot_input_router4) );
    AND2X1 U586 ( .IN1(new_rt_input_router4), .IN2(arst_valuenot_input_router4), .Q(finand3_input_router422) );
    MUX21X1 U587 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]), .IN2(next_rt_input_router4[0]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3]);
    MUX21X1 U588 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]), .IN2(next_rt_input_router4[1]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+1]);
    MUX21X1 U589 (.IN1(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]), .IN2(next_rt_input_router4[2]), .S(finand3_input_router422), .Q(routing_table_ff_input_router4[flit_input_router4_req_i[2]*3+2]); 


//input part


	BUFX1 U590 ( .A(read_ptr_ff_fifomodule[0]), .Y(next_read_ptr_fifomodule[0]) );
	BUFX1 U591 ( .A(read_ptr_ff_fifomodule[1]), .Y(next_read_ptr_fifomodule[1]) );
	BUFX1 U592 ( .A(write_ptr_ff_fifomodule[0]), .Y(next_write_ptr_fifomodule[0]) );
	BUFX1 U593 ( .A(write_ptr_ff_fifomodule[1]), .Y(next_write_ptr_fifomodule[1]) );

	XNOR2X1 U594 ( .IN1(write_ptr_ff_fifomodule[0]), .IN2(read_ptr_ff_fifomodule[0]), .Q(u1temp_fifomodule) );
	XNOR2X1 U595 ( .IN1(write_ptr_ff_fifomodule[1]), .IN2(read_ptr_ff_fifomodule[1]), .Q(u2temp_fifomodule) );
	AND2X1 U596 ( .A(u1temp_fifomodule), .B(u2temp_fifomodule), .Y(empty_vc_buffer) );
	XOR2X1 U597 ( .A(write_ptr_ff_fifomodule[1]), .B(read_ptr_ff_fifomodule[1]), .Y(u4temp_fifomodule) );
	AND2X1 U598 ( .A(u1temp_fifomodule), .B(u4temp_fifomodule), .Y(full_vc_buffer) );
	MUX21X1 U599 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][0]));
	MUX21X1 U600 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][1]));
	MUX21X1 U601 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][2]));
	MUX21X1 U602 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][3]));
	MUX21X1 U603 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][4]));
	MUX21X1 U604 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][5]));
	MUX21X1 U605 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][6]));
	MUX21X1 U606 (.IN1(fifo_ff_fifomodule[read_ptr_ff_fifomodule[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer), .Q(to_output_req_in_jump_input_datapathput_datapath[36:3][7]));

	INVX1 U607 ( .A(full_vc_buffer), .Y(full_vc_buffer_not_fifomodule) );
	AND2X1 U608 ( .A(write_flit_vc_buffer), .B(full_vc_buffer_not_fifomodule), .Y(u7temp_fifomodule) );
	MUX21X1 U609 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule), .Q(u9temp_fifomodule));
	HADDX1 U610 ( .A0(write_ptr_ff_fifomodule[0]), .B0(u9temp_fifomodule), .C1(u10carry_fifomodule), .SO(next_write_ptr_fifomodule[0]) );
	HADDX1 U611 ( .A0(u10carry_fifomodule), .B0(write_ptr_ff_fifomodule[1]), .C1(u11carry_fifomodule), .SO(next_write_ptr_fifomodule[1]) );

	INVX1 U612 ( .A(empty_vc_buffer), .Y(empty_vc_buffer_not_fifomodule) );
	AND2X1 U613 ( .A(read_flit_vc_buffer), .B(empty_vc_buffer_not_fifomodule), .Y(u13temp_fifomodule) );
	MUX21X1 U614 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule), .Q(u14temp_fifomodule));
	HADDX1 U615 ( .A0(read_ptr_ff_fifomodule[0]), .B0(u14temp_fifomodule), .C1(u15carry_fifomodule), .SO(next_read_ptr_fifomodule[0]) );
	HADDX1 U616 ( .A0(u15carry_fifomodule), .B0(read_ptr_ff_fifomodule[1]), .C1(u16carry_fifomodule), .SO(next_read_ptr_fifomodule[1]) );

	AND2X1 U617 ( .A(write_flit_vc_buffer), .B(full_vc_buffer), .Y(u17res_fifomodule) );
	AND2X1 U618 ( .A(read_flit_vc_buffer), .B(empty_vc_buffer), .Y(u18res_fifomodule) );
    OR2X1 U619 ( .A(u17res_fifomodule), .B(u18res_fifomodule), .Y(error_vc_buffer) );
	XOR2X1 U620 ( .A(write_ptr_ff_fifomodule[0]), .B(read_ptr_ff_fifomodule[0]), .Y(fifo_ocup_fifomodule[0]) );
	INVX1 U621 ( .A(write_ptr_ff_fifomodule[0]), .Y(write_ptr_ff_fifomodule_0_not) );
	AND2X1 U622 ( .A(write_ptr_ff_fifomodule_0_not), .B(read_ptr_ff_fifomodule[0]), .Y(b0wire_fifomodule) );
	XOR2X1 U623 ( .A(write_ptr_ff_fifomodule[1]), .B(read_ptr_ff_fifomodule[1]), .Y(u23temp_fifomodule) );
	INVX1 U624 ( .A(write_ptr_ff_fifomodule[1]), .Y(write_ptr_ff_fifomodule_1_not) );
	AND2X1 U625 ( .A(read_ptr_ff_fifomodule[1]), .B(write_ptr_ff_fifomodule_1_not), .Y(boutb_fifomodule) );
	XOR2X1 U626 ( .A(u23temp_fifomodule), .B(b0wire_fifomodule), .Y(fifo_ocup_fifomodule[1]) );
	INVX1 U627 ( .A(u23temp_fifomodule), .Y(u23temp_fifomodule_not_fifomodule) );
	AND2X1 U628 ( .A(b0wire_fifomodule), .B(u23temp_fifomodule_not_fifomodule), .Y(bouta_fifomodule) );
	OR2X1 U629 ( .A(bouta_fifomodule), .B(boutb_fifomodule), .Y(boutmain_fifomodule) );
	DFFX2 U630 ( .CLK(clk), .D(fifo_ocup_fifomodule[0]), .Q(ocup_o[0]) );
	DFFX2 U631 ( .CLK(clk), .D(fifo_ocup_fifomodule[1]), .Q(ocup_o[1]) );
	DFFX2 U632 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule) );
	DFFX2 U633 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule) );
	DFFX2 U634 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(write_ptr_ff_fifomodule[0]) );
	DFFX2 U635 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(read_ptr_ff_fifomodule[0]) );
	DFFX2 U636 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(fifo_ff_fifomodule[0]) );
	DFFX2 U637 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(write_ptr_ff_fifomodule[1]) );
	DFFX2 U638 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(read_ptr_ff_fifomodule[1]) );
	DFFX2 U639 ( .CLK(arst_value_fifomodule), .D(1'b0), .Q(fifo_ff_fifomodule[1]) );

	DFFX2 U640 ( .CLK(clk), .D(next_write_ptr_fifomodule[0]), .Q(write_ptr_ff_fifomodule[0]) );
	DFFX2 U641 ( .CLK(clk), .D(next_write_ptr_fifomodule[1]), .Q(write_ptr_ff_fifomodule[1]) );
	DFFX2 U642 ( .CLK(clk), .D(next_read_ptr_fifomodule[0]), .Q(read_ptr_ff_fifomodule[0]) );
	DFFX2 U643 ( .CLK(clk), .D(next_read_ptr_fifomodule[1]), .Q(read_ptr_ff_fifomodule[1]) );
	  

	DFFX2 U644 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][0]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8]) );
	DFFX2 U645 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][1]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+1]) );
	DFFX2 U646 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][2]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+2]) );
	DFFX2 U647 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][3]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+3]) );
	DFFX2 U648 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][4]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+4]) );
	DFFX2 U649 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][5]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+5]) );
	DFFX2 U650 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][6]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+6]) );
	DFFX2 U651 ( .CLK(u7temp_fifomodule), .D(from_input_req_in_jump_input_datapathput_datapath[36:3][7]), .Q(fifo_ff_fifomodule[write_ptr_ff_fifomodule[0]*8+7]) );

    BUFX1 U652 ( .A(locked_by_route_ff_vc_buffer), .Y(next_locked_vc_buffer) );
    BUFX1 U653(.A(flit[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][0]));
	BUFX1 U654(.A(flit[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][1]));
	BUFX1 U655(.A(flit[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][2]));
	BUFX1 U656(.A(flit[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][3]));
	BUFX1 U657(.A(flit[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][4]));
	BUFX1 U658(.A(flit[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][5]));
	BUFX1 U659(.A(flit[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][6]));
	BUFX1 U660(.A(flit[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][7]));
	BUFX1 U661(.A(flit[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][8]));
	BUFX1 U662(.A(flit[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][9]));
	BUFX1 U663(.A(flit[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][10]));
	BUFX1 U664(.A(flit[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][11]));
	BUFX1 U665(.A(flit[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][12]));
	BUFX1 U666(.A(flit[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][13]));
	BUFX1 U667(.A(flit[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][14]));
	BUFX1 U668(.A(flit[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][15]));
	BUFX1 U669(.A(flit[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][16]));
	BUFX1 U670(.A(flit[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][17]));
	BUFX1 U671(.A(flit[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][18]));
	BUFX1 U672(.A(flit[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][19]));
	BUFX1 U673(.A(flit[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][20]));
	BUFX1 U674(.A(flit[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][21]));
	BUFX1 U675(.A(flit[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][22]));
	BUFX1 U676(.A(flit[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][23]));
	BUFX1 U677(.A(flit[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][24]));
	BUFX1 U678(.A(flit[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][25]));
	BUFX1 U679(.A(flit[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][26]));
	BUFX1 U680(.A(flit[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][27]));
	BUFX1 U681(.A(flit[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][28]));
	BUFX1 U682(.A(flit[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][29]));
	BUFX1 U683(.A(flit[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][30]));
	BUFX1 U684(.A(flit[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][31]));
	BUFX1 U685(.A(flit[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][32]));
	BUFX1 U686(.A(flit[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[36:3][33]));
    NOR2X1 U687 ( .IN1(flit[33]), .IN2(flit[32]), .QN(norres_vc_buffer_vc_buffer) );
    OR4X1 U688 ( .IN1(flit[29]), .IN2(flit[28]), .IN3(flit[27]), .IN4(flit[26]), .Y(or1res_vc_buffer) );
    OR4X1 U689 ( .IN1(flit[25]), .IN2(flit[24]), .IN3(flit[23]), .IN4(flit[22]), .Y(or2res_vc_buffer) );
    OR2X1 U690 ( .A(or1res_vc_buffer), .B(or2res_vc_buffer), .Y(orres_vc_buffer) );
    AND3X1 U691 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(norres_vc_buffer_vc_buffer), .IN3(orres_vc_buffer), .Q(finres1_vc_buffer) );
    MUX21X1 U692 (.IN1(next_locked_vc_buffer), .IN2(1'b1), .S(finres1_vc_buffer), .Q(next_locked_vc_buffer);
    AND3X1 U693 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(flit[33]), .IN3(flit[32]), .Q(andres1_vc_buffer) );
    MUX21X1 U694 (.IN1(next_locked_vc_buffer), .IN2(1'b0), .S(andres1_vc_buffer), .Q(next_locked_vc_buffer);

    INVX1 U695 ( .A(full_vc_buffer), .Y(full_vc_buffer_not) );
    INVX1 U696 ( .A(locked_by_route_ff_vc_buffer), .Y(locked_by_route_ff_vc_buffer_not) );

    MUX21X1 U697 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer_not), .S(norres_vc_buffer_vc_buffer), .Q(thirdand_vc_buffer);
    AND3X1 U698 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[0]), .IN2(full_vc_buffer_not), .IN3(thirdand_vc_buffer), .Q(write_flit_vc_buffer) );
    AND2X1 U699 ( .IN1(full_vc_buffer_not), .IN2(norres_vc_buffer_vc_buffer), .Q(from_input_resp_input_datapath[0]) );
    INVX1 U700 ( .A(empty_vc_buffer), .Y(to_output_req_in_jump_input_datapathput_datapath[0]) );
    AND2X1 U701 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[0]), .IN2(to_output_resp_input_datapath[0]), .Q(read_flit_vc_buffer) );
	BUFX1 U702(.A(to_output_req_in_jump_input_datapathput_datapath[2:1]), .Y(2'b00));

	DFFX2 U703 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U704 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U705 (.IN1(next_locked_vc_buffer), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer);

	BUFX1 U706 ( .A(read_ptr_ff_fifomodule1[0]), .Y(next_read_ptr_fifomodule1[0]) );
	BUFX1 U707 ( .A(read_ptr_ff_fifomodule1[1]), .Y(next_read_ptr_fifomodule1[1]) );
	BUFX1 U708 ( .A(write_ptr_ff_fifomodule1[0]), .Y(next_write_ptr_fifomodule1[0]) );
	BUFX1 U709 ( .A(write_ptr_ff_fifomodule1[1]), .Y(next_write_ptr_fifomodule1[1]) );

	XNOR2X1 U710 ( .IN1(write_ptr_ff_fifomodule1[0]), .IN2(read_ptr_ff_fifomodule1[0]), .Q(u1temp_fifomodule1) );
	XNOR2X1 U711 ( .IN1(write_ptr_ff_fifomodule1[1]), .IN2(read_ptr_ff_fifomodule1[1]), .Q(u2temp_fifomodule1) );
	AND2X1 U712 ( .A(u1temp_fifomodule1), .B(u2temp_fifomodule1), .Y(empty_vc_buffer1) );
	XOR2X1 U713 ( .A(write_ptr_ff_fifomodule1[1]), .B(read_ptr_ff_fifomodule1[1]), .Y(u4temp_fifomodule1) );
	AND2X1 U714 ( .A(u1temp_fifomodule1), .B(u4temp_fifomodule1), .Y(full_vc_buffer1) );
	MUX21X1 U715 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][0]));
	MUX21X1 U716 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][1]));
	MUX21X1 U717 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][2]));
	MUX21X1 U718 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][3]));
	MUX21X1 U719 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][4]));
	MUX21X1 U720 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][5]));
	MUX21X1 U721 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][6]));
	MUX21X1 U722 (.IN1(fifo_ff_fifomodule1[read_ptr_ff_fifomodule1[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer1), .Q(to_output_req_in_jump_input_datapathput_datapath[73:40][7]));

	INVX1 U723 ( .A(full_vc_buffer1), .Y(full_vc_buffer1_not1_fifomodule1) );
	AND2X1 U724 ( .A(write_flit1_vc_buffer1), .B(full_vc_buffer1_not1_fifomodule1), .Y(u7temp_fifomodule1) );
	MUX21X1 U725 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule1), .Q(u9temp_fifomodule1));
	HADDX1 U726 ( .A0(write_ptr_ff_fifomodule1[0]), .B0(u9temp_fifomodule1), .C1(u10carry_fifomodule1), .SO(next_write_ptr_fifomodule1[0]) );
	HADDX1 U727 ( .A0(u10carry_fifomodule1), .B0(write_ptr_ff_fifomodule1[1]), .C1(u11carry_fifomodule1), .SO(next_write_ptr_fifomodule1[1]) );

	INVX1 U728 ( .A(empty_vc_buffer1), .Y(empty_vc_buffer1_not_fifomodule1) );
	AND2X1 U729 ( .A(read_flit1_vc_buffer1), .B(empty_vc_buffer1_not_fifomodule1), .Y(u13temp_fifomodule1) );
	MUX21X1 U730 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule1), .Q(u14temp_fifomodule1));
	HADDX1 U731 ( .A0(read_ptr_ff_fifomodule1[0]), .B0(u14temp_fifomodule1), .C1(u15carry_fifomodule1), .SO(next_read_ptr_fifomodule1[0]) );
	HADDX1 U732 ( .A0(u15carry_fifomodule1), .B0(read_ptr_ff_fifomodule1[1]), .C1(u16carry_fifomodule1), .SO(next_read_ptr_fifomodule1[1]) );

	AND2X1 U733 ( .A(write_flit1_vc_buffer1), .B(full_vc_buffer1), .Y(u17res_fifomodule1) );
	AND2X1 U734 ( .A(read_flit1_vc_buffer1), .B(empty_vc_buffer1), .Y(u18res_fifomodule1) );
    OR2X1 U735 ( .A(u17res_fifomodule1), .B(u18res_fifomodule1), .Y(error_vc_buffer1) );
	XOR2X1 U736 ( .A(write_ptr_ff_fifomodule1[0]), .B(read_ptr_ff_fifomodule1[0]), .Y(fifo_ocup_fifomodule1[0]) );
	INVX1 U737 ( .A(write_ptr_ff_fifomodule1[0]), .Y(write_ptr_ff_fifomodule1_0_not1) );
	AND2X1 U738 ( .A(write_ptr_ff_fifomodule1_0_not1), .B(read_ptr_ff_fifomodule1[0]), .Y(b0wire_fifomodule1) );
	XOR2X1 U739 ( .A(write_ptr_ff_fifomodule1[1]), .B(read_ptr_ff_fifomodule1[1]), .Y(u23temp_fifomodule1) );
	INVX1 U740 ( .A(write_ptr_ff_fifomodule1[1]), .Y(write_ptr_ff_fifomodule1_1_not1) );
	AND2X1 U741 ( .A(read_ptr_ff_fifomodule1[1]), .B(write_ptr_ff_fifomodule1_1_not1), .Y(boutb_fifomodule1) );
	XOR2X1 U742 ( .A(u23temp_fifomodule1), .B(b0wire_fifomodule1), .Y(fifo_ocup_fifomodule1[1]) );
	INVX1 U743 ( .A(u23temp_fifomodule1), .Y(u23temp_fifomodule1_not_fifomodule1) );
	AND2X1 U744 ( .A(b0wire_fifomodule1), .B(u23temp_fifomodule1_not_fifomodule1), .Y(bouta_fifomodule1) );
	OR2X1 U745 ( .A(bouta_fifomodule1), .B(boutb_fifomodule1), .Y(boutmain_fifomodule1) );
	DFFX2 U746 ( .CLK(clk), .D(fifo_ocup_fifomodule1[0]), .Q(ocup_o[0]) );
	DFFX2 U747 ( .CLK(clk), .D(fifo_ocup_fifomodule1[1]), .Q(ocup_o[1]) );
	DFFX2 U748 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule1) );
	DFFX2 U749 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule1) );
	DFFX2 U750 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(write_ptr_ff_fifomodule1[0]) );
	DFFX2 U751 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(read_ptr_ff_fifomodule1[0]) );
	DFFX2 U752 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(fifo_ff_fifomodule1[0]) );
	DFFX2 U753 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(write_ptr_ff_fifomodule1[1]) );
	DFFX2 U754 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(read_ptr_ff_fifomodule1[1]) );
	DFFX2 U755 ( .CLK(arst_value_fifomodule1), .D(1'b0), .Q(fifo_ff_fifomodule1[1]) );

	DFFX2 U756 ( .CLK(clk), .D(next_write_ptr_fifomodule1[0]), .Q(write_ptr_ff_fifomodule1[0]) );
	DFFX2 U757 ( .CLK(clk), .D(next_write_ptr_fifomodule1[1]), .Q(write_ptr_ff_fifomodule1[1]) );
	DFFX2 U758 ( .CLK(clk), .D(next_read_ptr_fifomodule1[0]), .Q(read_ptr_ff_fifomodule1[0]) );
	DFFX2 U759 ( .CLK(clk), .D(next_read_ptr_fifomodule1[1]), .Q(read_ptr_ff_fifomodule1[1]) );
	  

	DFFX2 U760 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][0]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8]) );
	DFFX2 U761 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][1]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+1]) );
	DFFX2 U762 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][2]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+2]) );
	DFFX2 U763 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][3]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+3]) );
	DFFX2 U764 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][4]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+4]) );
	DFFX2 U765 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][5]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+5]) );
	DFFX2 U766 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][6]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+6]) );
	DFFX2 U767 ( .CLK(u7temp_fifomodule1), .D(from_input_req_in_jump_input_datapathput_datapath[73:40][7]), .Q(fifo_ff_fifomodule1[write_ptr_ff_fifomodule1[0]*8+7]) );

    BUFX1 U768 ( .A(locked_by_route_ff_vc_buffer1), .Y(next_locked_vc_buffer1) );
    BUFX1 U769(.A(flit1[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][0]));
	BUFX1 U770(.A(flit1[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][1]));
	BUFX1 U771(.A(flit1[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][2]));
	BUFX1 U772(.A(flit1[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][3]));
	BUFX1 U773(.A(flit1[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][4]));
	BUFX1 U774(.A(flit1[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][5]));
	BUFX1 U775(.A(flit1[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][6]));
	BUFX1 U776(.A(flit1[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][7]));
	BUFX1 U777(.A(flit1[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][8]));
	BUFX1 U778(.A(flit1[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][9]));
	BUFX1 U779(.A(flit1[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][10]));
	BUFX1 U780(.A(flit1[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][11]));
	BUFX1 U781(.A(flit1[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][12]));
	BUFX1 U782(.A(flit1[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][13]));
	BUFX1 U783(.A(flit1[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][14]));
	BUFX1 U784(.A(flit1[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][15]));
	BUFX1 U785(.A(flit1[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][16]));
	BUFX1 U786(.A(flit1[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][17]));
	BUFX1 U787(.A(flit1[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][18]));
	BUFX1 U788(.A(flit1[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][19]));
	BUFX1 U789(.A(flit1[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][20]));
	BUFX1 U790(.A(flit1[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][21]));
	BUFX1 U791(.A(flit1[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][22]));
	BUFX1 U792(.A(flit1[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][23]));
	BUFX1 U793(.A(flit1[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][24]));
	BUFX1 U794(.A(flit1[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][25]));
	BUFX1 U795(.A(flit1[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][26]));
	BUFX1 U796(.A(flit1[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][27]));
	BUFX1 U797(.A(flit1[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][28]));
	BUFX1 U798(.A(flit1[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][29]));
	BUFX1 U799(.A(flit1[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][30]));
	BUFX1 U800(.A(flit1[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][31]));
	BUFX1 U801(.A(flit1[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][32]));
	BUFX1 U802(.A(flit1[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[73:40][33]));
    NOR2X1 U803 ( .IN1(flit1[33]), .IN2(flit1[32]), .QN(norres_vc_buffer1_vc_buffer1) );
    OR4X1 U804 ( .IN1(flit1[29]), .IN2(flit1[28]), .IN3(flit1[27]), .IN4(flit1[26]), .Y(or1res_vc_buffer1) );
    OR4X1 U805 ( .IN1(flit1[25]), .IN2(flit1[24]), .IN3(flit1[23]), .IN4(flit1[22]), .Y(or2res_vc_buffer1) );
    OR2X1 U806 ( .A(or1res_vc_buffer1), .B(or2res_vc_buffer1), .Y(orres_vc_buffer1) );
    AND3X1 U807 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(norres_vc_buffer1_vc_buffer1), .IN3(orres_vc_buffer1), .Q(finres1_vc_buffer1) );
    MUX21X1 U808 (.IN1(next_locked_vc_buffer1), .IN2(1'b1), .S(finres1_vc_buffer1), .Q(next_locked_vc_buffer1);
    AND3X1 U809 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(flit1[33]), .IN3(flit1[32]), .Q(andres1_vc_buffer1) );
    MUX21X1 U810 (.IN1(next_locked_vc_buffer1), .IN2(1'b0), .S(andres1_vc_buffer1), .Q(next_locked_vc_buffer1);

    INVX1 U811 ( .A(full_vc_buffer1), .Y(full_vc_buffer1_not1) );
    INVX1 U812 ( .A(locked_by_route_ff_vc_buffer1), .Y(locked_by_route_ff_vc_buffer1_not1) );

    MUX21X1 U813 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer1_not1), .S(norres_vc_buffer1_vc_buffer1), .Q(thirdand_vc_buffer1);
    AND3X1 U814 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[37]), .IN2(full_vc_buffer1_not1), .IN3(thirdand_vc_buffer1), .Q(write_flit1_vc_buffer1) );
    AND2X1 U815 ( .IN1(full_vc_buffer1_not1), .IN2(norres_vc_buffer1_vc_buffer1), .Q(from_input_resp_input_datapath[1]) );
    INVX1 U816 ( .A(empty_vc_buffer1), .Y(to_output_req_in_jump_input_datapathput_datapath[37]) );
    AND2X1 U817 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[37]), .IN2(to_output_resp_input_datapath[1]), .Q(read_flit1_vc_buffer1) );
	BUFX1 U818(.A(to_output_req_in_jump_input_datapathput_datapath[39:38]), .Y(2'b01));

	DFFX2 U819 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U820 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U821 (.IN1(next_locked_vc_buffer1), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer1);


	BUFX1 U822 ( .A(read_ptr_ff_fifomodule2[0]), .Y(next_read_ptr_fifomodule2[0]) );
	BUFX1 U823 ( .A(read_ptr_ff_fifomodule2[1]), .Y(next_read_ptr_fifomodule2[1]) );
	BUFX1 U824 ( .A(write_ptr_ff_fifomodule2[0]), .Y(next_write_ptr_fifomodule2[0]) );
	BUFX1 U825 ( .A(write_ptr_ff_fifomodule2[1]), .Y(next_write_ptr_fifomodule2[1]) );

	XNOR2X1 U826 ( .IN1(write_ptr_ff_fifomodule2[0]), .IN2(read_ptr_ff_fifomodule2[0]), .Q(u1temp_fifomodule2) );
	XNOR2X1 U827 ( .IN1(write_ptr_ff_fifomodule2[1]), .IN2(read_ptr_ff_fifomodule2[1]), .Q(u2temp_fifomodule2) );
	AND2X1 U828 ( .A(u1temp_fifomodule2), .B(u2temp_fifomodule2), .Y(empty_vc_buffer2) );
	XOR2X1 U829 ( .A(write_ptr_ff_fifomodule2[1]), .B(read_ptr_ff_fifomodule2[1]), .Y(u4temp_fifomodule2) );
	AND2X1 U830 ( .A(u1temp_fifomodule2), .B(u4temp_fifomodule2), .Y(full_vc_buffer2) );
	MUX21X1 U831 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][0]));
	MUX21X1 U832 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][1]));
	MUX21X1 U833 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][2]));
	MUX21X1 U834 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][3]));
	MUX21X1 U835 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][4]));
	MUX21X1 U836 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][5]));
	MUX21X1 U837 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][6]));
	MUX21X1 U838 (.IN1(fifo_ff_fifomodule2[read_ptr_ff_fifomodule2[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer2), .Q(to_output_req_in_jump_input_datapathput_datapath[110:77][7]));

	INVX1 U839 ( .A(full_vc_buffer2), .Y(full_vc_buffer2_not2_fifomodule2) );
	AND2X1 U840 ( .A(write_flit2_vc_buffer2), .B(full_vc_buffer2_not2_fifomodule2), .Y(u7temp_fifomodule2) );
	MUX21X1 U841 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule2), .Q(u9temp_fifomodule2));
	HADDX1 U842 ( .A0(write_ptr_ff_fifomodule2[0]), .B0(u9temp_fifomodule2), .C1(u10carry_fifomodule2), .SO(next_write_ptr_fifomodule2[0]) );
	HADDX1 U843 ( .A0(u10carry_fifomodule2), .B0(write_ptr_ff_fifomodule2[1]), .C1(u11carry_fifomodule2), .SO(next_write_ptr_fifomodule2[1]) );

	INVX1 U844 ( .A(empty_vc_buffer2), .Y(empty_vc_buffer2_not_fifomodule2) );
	AND2X1 U845 ( .A(read_flit2_vc_buffer2), .B(empty_vc_buffer2_not_fifomodule2), .Y(u13temp_fifomodule2) );
	MUX21X1 U846 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule2), .Q(u14temp_fifomodule2));
	HADDX1 U847 ( .A0(read_ptr_ff_fifomodule2[0]), .B0(u14temp_fifomodule2), .C1(u15carry_fifomodule2), .SO(next_read_ptr_fifomodule2[0]) );
	HADDX1 U848 ( .A0(u15carry_fifomodule2), .B0(read_ptr_ff_fifomodule2[1]), .C1(u16carry_fifomodule2), .SO(next_read_ptr_fifomodule2[1]) );

	AND2X1 U849 ( .A(write_flit2_vc_buffer2), .B(full_vc_buffer2), .Y(u17res_fifomodule2) );
	AND2X1 U850 ( .A(read_flit2_vc_buffer2), .B(empty_vc_buffer2), .Y(u18res_fifomodule2) );
    OR2X1 U851 ( .A(u17res_fifomodule2), .B(u18res_fifomodule2), .Y(error_vc_buffer2) );
	XOR2X1 U852 ( .A(write_ptr_ff_fifomodule2[0]), .B(read_ptr_ff_fifomodule2[0]), .Y(fifo_ocup_fifomodule2[0]) );
	INVX1 U853 ( .A(write_ptr_ff_fifomodule2[0]), .Y(write_ptr_ff_fifomodule2_0_not2) );
	AND2X1 U854 ( .A(write_ptr_ff_fifomodule2_0_not2), .B(read_ptr_ff_fifomodule2[0]), .Y(b0wire_fifomodule2) );
	XOR2X1 U855 ( .A(write_ptr_ff_fifomodule2[1]), .B(read_ptr_ff_fifomodule2[1]), .Y(u23temp_fifomodule2) );
	INVX1 U856 ( .A(write_ptr_ff_fifomodule2[1]), .Y(write_ptr_ff_fifomodule2_1_not2) );
	AND2X1 U857 ( .A(read_ptr_ff_fifomodule2[1]), .B(write_ptr_ff_fifomodule2_1_not2), .Y(boutb_fifomodule2) );
	XOR2X1 U858 ( .A(u23temp_fifomodule2), .B(b0wire_fifomodule2), .Y(fifo_ocup_fifomodule2[1]) );
	INVX1 U859 ( .A(u23temp_fifomodule2), .Y(u23temp_fifomodule2_not_fifomodule2) );
	AND2X1 U860 ( .A(b0wire_fifomodule2), .B(u23temp_fifomodule2_not_fifomodule2), .Y(bouta_fifomodule2) );
	OR2X1 U861 ( .A(bouta_fifomodule2), .B(boutb_fifomodule2), .Y(boutmain_fifomodule2) );
	DFFX2 U862 ( .CLK(clk), .D(fifo_ocup_fifomodule2[0]), .Q(ocup_o[0]) );
	DFFX2 U863 ( .CLK(clk), .D(fifo_ocup_fifomodule2[1]), .Q(ocup_o[1]) );
	DFFX2 U864 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule2) );
	DFFX2 U865 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule2) );
	DFFX2 U866 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(write_ptr_ff_fifomodule2[0]) );
	DFFX2 U867 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(read_ptr_ff_fifomodule2[0]) );
	DFFX2 U868 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(fifo_ff_fifomodule2[0]) );
	DFFX2 U869 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(write_ptr_ff_fifomodule2[1]) );
	DFFX2 U870 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(read_ptr_ff_fifomodule2[1]) );
	DFFX2 U871 ( .CLK(arst_value_fifomodule2), .D(1'b0), .Q(fifo_ff_fifomodule2[1]) );

	DFFX2 U872 ( .CLK(clk), .D(next_write_ptr_fifomodule2[0]), .Q(write_ptr_ff_fifomodule2[0]) );
	DFFX2 U873 ( .CLK(clk), .D(next_write_ptr_fifomodule2[1]), .Q(write_ptr_ff_fifomodule2[1]) );
	DFFX2 U874 ( .CLK(clk), .D(next_read_ptr_fifomodule2[0]), .Q(read_ptr_ff_fifomodule2[0]) );
	DFFX2 U875 ( .CLK(clk), .D(next_read_ptr_fifomodule2[1]), .Q(read_ptr_ff_fifomodule2[1]) );
	  

	DFFX2 U876 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][0]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8]) );
	DFFX2 U877 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][1]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+1]) );
	DFFX2 U878 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][2]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+2]) );
	DFFX2 U879 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][3]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+3]) );
	DFFX2 U880 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][4]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+4]) );
	DFFX2 U881 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][5]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+5]) );
	DFFX2 U882 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][6]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+6]) );
	DFFX2 U883 ( .CLK(u7temp_fifomodule2), .D(from_input_req_in_jump_input_datapathput_datapath[110:77][7]), .Q(fifo_ff_fifomodule2[write_ptr_ff_fifomodule2[0]*8+7]) );

    BUFX1 U884 ( .A(locked_by_route_ff_vc_buffer2), .Y(next_locked_vc_buffer2) );
    BUFX1 U885(.A(flit2[0]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][0]));
	BUFX1 U886(.A(flit2[1]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][1]));
	BUFX1 U887(.A(flit2[2]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][2]));
	BUFX1 U888(.A(flit2[3]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][3]));
	BUFX1 U889(.A(flit2[4]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][4]));
	BUFX1 U890(.A(flit2[5]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][5]));
	BUFX1 U891(.A(flit2[6]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][6]));
	BUFX1 U892(.A(flit2[7]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][7]));
	BUFX1 U893(.A(flit2[8]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][8]));
	BUFX1 U894(.A(flit2[9]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][9]));
	BUFX1 U895(.A(flit2[10]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][10]));
	BUFX1 U896(.A(flit2[11]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][11]));
	BUFX1 U897(.A(flit2[12]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][12]));
	BUFX1 U898(.A(flit2[13]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][13]));
	BUFX1 U899(.A(flit2[14]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][14]));
	BUFX1 U900(.A(flit2[15]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][15]));
	BUFX1 U901(.A(flit2[16]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][16]));
	BUFX1 U902(.A(flit2[17]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][17]));
	BUFX1 U903(.A(flit2[18]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][18]));
	BUFX1 U904(.A(flit2[19]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][19]));
	BUFX1 U905(.A(flit2[20]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][20]));
	BUFX1 U906(.A(flit2[21]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][21]));
	BUFX1 U907(.A(flit2[22]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][22]));
	BUFX1 U908(.A(flit2[23]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][23]));
	BUFX1 U909(.A(flit2[24]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][24]));
	BUFX1 U910(.A(flit2[25]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][25]));
	BUFX1 U911(.A(flit2[26]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][26]));
	BUFX1 U912(.A(flit2[27]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][27]));
	BUFX1 U913(.A(flit2[28]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][28]));
	BUFX1 U914(.A(flit2[29]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][29]));
	BUFX1 U915(.A(flit2[30]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][30]));
	BUFX1 U916(.A(flit2[31]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][31]));
	BUFX1 U917(.A(flit2[32]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][32]));
	BUFX1 U918(.A(flit2[33]), .Y(from_input_req_in_jump_input_datapathput_datapath[110:77][33]));
    NOR2X1 U919 ( .IN1(flit2[33]), .IN2(flit2[32]), .QN(norres_vc_buffer2_vc_buffer2) );
    OR4X1 U920 ( .IN1(flit2[29]), .IN2(flit2[28]), .IN3(flit2[27]), .IN4(flit2[26]), .Y(or1res_vc_buffer2) );
    OR4X1 U921 ( .IN1(flit2[25]), .IN2(flit2[24]), .IN3(flit2[23]), .IN4(flit2[22]), .Y(or2res_vc_buffer2) );
    OR2X1 U922 ( .A(or1res_vc_buffer2), .B(or2res_vc_buffer2), .Y(orres_vc_buffer2) );
    AND3X1 U923 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(norres_vc_buffer2_vc_buffer2), .IN3(orres_vc_buffer2), .Q(finres1_vc_buffer2) );
    MUX21X1 U924 (.IN1(next_locked_vc_buffer2), .IN2(1'b1), .S(finres1_vc_buffer2), .Q(next_locked_vc_buffer2);
    AND3X1 U925 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(flit2[33]), .IN3(flit2[32]), .Q(andres1_vc_buffer2) );
    MUX21X1 U926 (.IN1(next_locked_vc_buffer2), .IN2(1'b0), .S(andres1_vc_buffer2), .Q(next_locked_vc_buffer2);

    INVX1 U927 ( .A(full_vc_buffer2), .Y(full_vc_buffer2_not2) );
    INVX1 U928 ( .A(locked_by_route_ff_vc_buffer2), .Y(locked_by_route_ff_vc_buffer2_not2) );

    MUX21X1 U929 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer2_not2), .S(norres_vc_buffer2_vc_buffer2), .Q(thirdand_vc_buffer2);
    AND3X1 U930 ( .IN1(from_input_req_in_jump_input_datapathput_datapath[74]), .IN2(full_vc_buffer2_not2), .IN3(thirdand_vc_buffer2), .Q(write_flit2_vc_buffer2) );
    AND2X1 U931 ( .IN1(full_vc_buffer2_not2), .IN2(norres_vc_buffer2_vc_buffer2), .Q(from_input_resp_input_datapath[2]) );
    INVX1 U932 ( .A(empty_vc_buffer2), .Y(to_output_req_in_jump_input_datapathput_datapath[74]) );
    AND2X1 U933 ( .IN1(to_output_req_in_jump_input_datapathput_datapath[74]), .IN2(to_output_resp_input_datapath[2]), .Q(read_flit2_vc_buffer2) );
	BUFX1 U934(.A(to_output_req_in_jump_input_datapathput_datapath[76:75]), .Y(2'b10));

	DFFX2 U935 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U936 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U937 (.IN1(next_locked_vc_buffer2), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer2);

	BUFX1 U938(.A(from_input_req_in_jump_input_datapathput_datapath[77]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U939(.A(from_input_req_in_jump_input_datapathput_datapath[78]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U940(.A(from_input_req_in_jump_input_datapathput_datapath[79]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U941(.A(from_input_req_in_jump_input_datapathput_datapath[80]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U942(.A(from_input_req_in_jump_input_datapathput_datapath[81]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U943(.A(from_input_req_in_jump_input_datapathput_datapath[82]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U944(.A(from_input_req_in_jump_input_datapathput_datapath[83]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U945(.A(from_input_req_in_jump_input_datapathput_datapath[84]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U946(.A(from_input_req_in_jump_input_datapathput_datapath[85]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U947(.A(from_input_req_in_jump_input_datapathput_datapath[86]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U948(.A(from_input_req_in_jump_input_datapathput_datapath[87]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U949(.A(from_input_req_in_jump_input_datapathput_datapath[88]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U950(.A(from_input_req_in_jump_input_datapathput_datapath[89]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U951(.A(from_input_req_in_jump_input_datapathput_datapath[90]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U952(.A(from_input_req_in_jump_input_datapathput_datapath[91]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U953(.A(from_input_req_in_jump_input_datapathput_datapath[92]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U954(.A(from_input_req_in_jump_input_datapathput_datapath[93]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U955(.A(from_input_req_in_jump_input_datapathput_datapath[94]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U956(.A(from_input_req_in_jump_input_datapathput_datapath[95]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U957(.A(from_input_req_in_jump_input_datapathput_datapath[96]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U958(.A(from_input_req_in_jump_input_datapathput_datapath[97]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U959(.A(from_input_req_in_jump_input_datapathput_datapath[98]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U960(.A(from_input_req_in_jump_input_datapathput_datapath[99]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U961(.A(from_input_req_in_jump_input_datapathput_datapath[100]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U962(.A(from_input_req_in_jump_input_datapathput_datapath[101]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U963(.A(from_input_req_in_jump_input_datapathput_datapath[102]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U964(.A(from_input_req_in_jump_input_datapathput_datapath[103]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U965(.A(from_input_req_in_jump_input_datapathput_datapath[104]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U966(.A(from_input_req_in_jump_input_datapathput_datapath[105]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U967(.A(from_input_req_in_jump_input_datapathput_datapath[106]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U968(.A(from_input_req_in_jump_input_datapathput_datapath[107]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U969(.A(from_input_req_in_jump_input_datapathput_datapath[108]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U970(.A(from_input_req_in_jump_input_datapathput_datapath[109]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U971(.A(from_input_req_in_jump_input_datapathput_datapath[110]), .Y(ext_req_v_i[36:0][36]));
    XNOR2X1 U972 ( .IN1(ext_req_v_i[36:0][1]), .IN2(i_input_datapath[0]), .QN(xnor1resu_input_datapath) );
    XNOR2X1 U973 ( .IN1(ext_req_v_i[36:0][2]), .IN2(i_input_datapath[1]), .QN(xnor2resu_input_datapath) );
    AND2X1 U974 ( .IN1(xnor1resu_input_datapath), .IN2(xnor2resu_input_datapath), .Q(and1resu_input_datapath) );
    AND3X1 U975 ( .IN1(and1resu_input_datapath), .IN2(ext_req_v_i[36:0][0]), .IN2(ext_req_v_i[36:0][0]), .Q(cond1line_input_datapath) );
    MUX21X1 U976 (.IN1(vc_ch_act_in_input_datapath[0]), .IN2(i_input_datapath[0]), .S(cond1line_input_datapath), .Q(vc_ch_act_in_input_datapath[0]));
    MUX21X1 U977 (.IN1(vc_ch_act_in_input_datapath[1]), .IN2(i_input_datapath[1]), .S(cond1line_input_datapath), .Q(vc_ch_act_in_input_datapath[1]));
    MUX21X1 U978 (.IN1(req_in_jump_input_datapath), .IN2(1), .S(cond1line_input_datapath), .Q(req_in_jump_input_datapath));
	BUFX1 U979(.A(from_input_req_in_jump_input_datapathput_datapath[40]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U980(.A(from_input_req_in_jump_input_datapathput_datapath[41]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U981(.A(from_input_req_in_jump_input_datapathput_datapath[42]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U982(.A(from_input_req_in_jump_input_datapathput_datapath[43]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U983(.A(from_input_req_in_jump_input_datapathput_datapath[44]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U984(.A(from_input_req_in_jump_input_datapathput_datapath[45]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U985(.A(from_input_req_in_jump_input_datapathput_datapath[46]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U986(.A(from_input_req_in_jump_input_datapathput_datapath[47]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U987(.A(from_input_req_in_jump_input_datapathput_datapath[48]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U988(.A(from_input_req_in_jump_input_datapathput_datapath[49]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U989(.A(from_input_req_in_jump_input_datapathput_datapath[50]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U990(.A(from_input_req_in_jump_input_datapathput_datapath[51]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U991(.A(from_input_req_in_jump_input_datapathput_datapath[52]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U992(.A(from_input_req_in_jump_input_datapathput_datapath[53]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U993(.A(from_input_req_in_jump_input_datapathput_datapath[54]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U994(.A(from_input_req_in_jump_input_datapathput_datapath[55]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U995(.A(from_input_req_in_jump_input_datapathput_datapath[56]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U996(.A(from_input_req_in_jump_input_datapathput_datapath[57]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U997(.A(from_input_req_in_jump_input_datapathput_datapath[58]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U998(.A(from_input_req_in_jump_input_datapathput_datapath[59]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U999(.A(from_input_req_in_jump_input_datapathput_datapath[60]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U1000(.A(from_input_req_in_jump_input_datapathput_datapath[61]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U1001(.A(from_input_req_in_jump_input_datapathput_datapath[62]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U1002(.A(from_input_req_in_jump_input_datapathput_datapath[63]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U1003(.A(from_input_req_in_jump_input_datapathput_datapath[64]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U1004(.A(from_input_req_in_jump_input_datapathput_datapath[65]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U1005(.A(from_input_req_in_jump_input_datapathput_datapath[66]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U1006(.A(from_input_req_in_jump_input_datapathput_datapath[67]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U1007(.A(from_input_req_in_jump_input_datapathput_datapath[68]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U1008(.A(from_input_req_in_jump_input_datapathput_datapath[69]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U1009(.A(from_input_req_in_jump_input_datapathput_datapath[70]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U1010(.A(from_input_req_in_jump_input_datapathput_datapath[71]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U1011(.A(from_input_req_in_jump_input_datapathput_datapath[72]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U1012(.A(from_input_req_in_jump_input_datapathput_datapath[73]), .Y(ext_req_v_i[36:0][36]));

	BUFX1 U1013(.A(from_input_req_in_jump_input_datapathput_datapath[3]), .Y(ext_req_v_i[36:0][3]));
	BUFX1 U1014(.A(from_input_req_in_jump_input_datapathput_datapath[4]), .Y(ext_req_v_i[36:0][4]));
	BUFX1 U1015(.A(from_input_req_in_jump_input_datapathput_datapath[5]), .Y(ext_req_v_i[36:0][5]));
	BUFX1 U1016(.A(from_input_req_in_jump_input_datapathput_datapath[6]), .Y(ext_req_v_i[36:0][6]));
	BUFX1 U1017(.A(from_input_req_in_jump_input_datapathput_datapath[7]), .Y(ext_req_v_i[36:0][7]));
	BUFX1 U1018(.A(from_input_req_in_jump_input_datapathput_datapath[8]), .Y(ext_req_v_i[36:0][8]));
	BUFX1 U1019(.A(from_input_req_in_jump_input_datapathput_datapath[9]), .Y(ext_req_v_i[36:0][9]));
	BUFX1 U1020(.A(from_input_req_in_jump_input_datapathput_datapath[10]), .Y(ext_req_v_i[36:0][10]));
	BUFX1 U1021(.A(from_input_req_in_jump_input_datapathput_datapath[11]), .Y(ext_req_v_i[36:0][11]));
	BUFX1 U1022(.A(from_input_req_in_jump_input_datapathput_datapath[12]), .Y(ext_req_v_i[36:0][12]));
	BUFX1 U1023(.A(from_input_req_in_jump_input_datapathput_datapath[13]), .Y(ext_req_v_i[36:0][13]));
	BUFX1 U1024(.A(from_input_req_in_jump_input_datapathput_datapath[14]), .Y(ext_req_v_i[36:0][14]));
	BUFX1 U1025(.A(from_input_req_in_jump_input_datapathput_datapath[15]), .Y(ext_req_v_i[36:0][15]));
	BUFX1 U1026(.A(from_input_req_in_jump_input_datapathput_datapath[16]), .Y(ext_req_v_i[36:0][16]));
	BUFX1 U1027(.A(from_input_req_in_jump_input_datapathput_datapath[17]), .Y(ext_req_v_i[36:0][17]));
	BUFX1 U1028(.A(from_input_req_in_jump_input_datapathput_datapath[18]), .Y(ext_req_v_i[36:0][18]));
	BUFX1 U1029(.A(from_input_req_in_jump_input_datapathput_datapath[19]), .Y(ext_req_v_i[36:0][19]));
	BUFX1 U1030(.A(from_input_req_in_jump_input_datapathput_datapath[20]), .Y(ext_req_v_i[36:0][20]));
	BUFX1 U1031(.A(from_input_req_in_jump_input_datapathput_datapath[21]), .Y(ext_req_v_i[36:0][21]));
	BUFX1 U1032(.A(from_input_req_in_jump_input_datapathput_datapath[22]), .Y(ext_req_v_i[36:0][22]));
	BUFX1 U1033(.A(from_input_req_in_jump_input_datapathput_datapath[23]), .Y(ext_req_v_i[36:0][23]));
	BUFX1 U1034(.A(from_input_req_in_jump_input_datapathput_datapath[24]), .Y(ext_req_v_i[36:0][24]));
	BUFX1 U1035(.A(from_input_req_in_jump_input_datapathput_datapath[25]), .Y(ext_req_v_i[36:0][25]));
	BUFX1 U1036(.A(from_input_req_in_jump_input_datapathput_datapath[26]), .Y(ext_req_v_i[36:0][26]));
	BUFX1 U1037(.A(from_input_req_in_jump_input_datapathput_datapath[27]), .Y(ext_req_v_i[36:0][27]));
	BUFX1 U1038(.A(from_input_req_in_jump_input_datapathput_datapath[28]), .Y(ext_req_v_i[36:0][28]));
	BUFX1 U1039(.A(from_input_req_in_jump_input_datapathput_datapath[29]), .Y(ext_req_v_i[36:0][29]));
	BUFX1 U1040(.A(from_input_req_in_jump_input_datapathput_datapath[30]), .Y(ext_req_v_i[36:0][30]));
	BUFX1 U1041(.A(from_input_req_in_jump_input_datapathput_datapath[31]), .Y(ext_req_v_i[36:0][31]));
	BUFX1 U1042(.A(from_input_req_in_jump_input_datapathput_datapath[32]), .Y(ext_req_v_i[36:0][32]));
	BUFX1 U1043(.A(from_input_req_in_jump_input_datapathput_datapath[33]), .Y(ext_req_v_i[36:0][33]));
	BUFX1 U1044(.A(from_input_req_in_jump_input_datapathput_datapath[34]), .Y(ext_req_v_i[36:0][34]));
	BUFX1 U1045(.A(from_input_req_in_jump_input_datapathput_datapath[35]), .Y(ext_req_v_i[36:0][35]));
	BUFX1 U1046(.A(from_input_req_in_jump_input_datapathput_datapath[36]), .Y(ext_req_v_i[36:0][36]));

    MUX21X1 U1047 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath * 37]), .IN2(ext_req_v_i[36:0][0]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath * 37]));
    MUX21X1 U1048 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+2]), .IN2(vc_ch_act_in_input_datapath[1]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+2]));
    MUX21X1 U1049 (.IN1(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+1]), .IN2(vc_ch_act_in_input_datapath[0]), .S(req_in_jump_input_datapath), .Q(from_input_req_in_jump_input_datapathput_datapath[vc_ch_act_in_input_datapath*37+1]));
    MUX21X1 U1050 (.IN1(ext_resp_v_o[1:0][0]), .IN2(from_input_resp_input_datapath[vc_ch_act_in_input_datapath]), .S(req_in_jump_input_datapath), .Q(ext_resp_v_o[1:0][0]));

    INVX1 U1051 ( .A(req_in_jump_input_datapath), .Y(req_in_jump_input_datapath_not) );
    MUX21X1 U1052 (.IN1(ext_resp_v_o[1:0][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath_not), .Q(ext_resp_v_o[1:0][0]));
    BUFX1 U1053(.A(from_input_req_in_jump_input_datapathput_datapath[34]), .Y(ext_req_v_i[36:0][34]));

    XOR2X1 U1054 ( .IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b1), .Q(xor1resu_input_datapath) );
    MUX21X1 U1055 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(xor1resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U1056 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b0), .S(xor1resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    AND2X1 U1057 ( .IN1(xor1resu_input_datapath), .IN2(to_output_req_in_jump_input_datapathput_datapath[j_input_datapath*37]), .Q(and2resu_input_datapath) );
    MUX21X1 U1058 (.IN1(vc_ch_act_out_input_datapath[0]), .IN2(j_input_datapath[0]), .S(and2resu_input_datapath), .Q(vc_ch_act_out_input_datapath[0]));
    MUX21X1 U1059 (.IN1(vc_ch_act_out_input_datapath[1]), .IN2(j_input_datapath[1]), .S(and2resu_input_datapath), .Q(vc_ch_act_out_input_datapath[1]));
    MUX21X1 U1060 (.IN1(req_out_jump_input_datapath), .IN2(1'b1), .S(and2resu_input_datapath), .Q(req_out_jump_input_datapath));
    MUX21X1 U1061 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(and2resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U1062 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b1), .S(and2resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    HADDX1 U1063 ( .A0(j_input_datapath[0]), .B0(1'b1), .C1(j_input_datapath[1]), .SO(j_input_datapath[0]) );
    HADDX1 U1064 ( .A0(j_input_datapath[0]), .B0(1'b1), .C1(j_input_datapath[1]), .SO(j_input_datapath[0]) );
    AND2X1 U1065 ( .IN1(xor1resu_input_datapath), .IN2(to_output_req_in_jump_input_datapathput_datapath[j_input_datapath*37]), .Q(and3resu) );
    NAND2X1 U1066(.A(_sv2v_jump_input_datapath[0]),.B(_sv2v_jump_input_datapath[1]),.Y(nand1resu_input_datapath));
    MUX21X1 U1067 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(1'b0), .S(nand1resu_input_datapath), .Q(_sv2v_jump_input_datapath[0]));
    MUX21X1 U1068 (.IN1(_sv2v_jump_input_datapath[1]), .IN2(1'b0), .S(nand1resu_input_datapath), .Q(_sv2v_jump_input_datapath[1]));
    XNOR2X1 U1069 (.IN1(_sv2v_jump_input_datapath[0]), .IN2(_sv2v_jump_input_datapath[1]), .Q(xnor23resu_input_datapath) );
    AND2X1 U1070 ( .IN1(xnor23resu_input_datapath), .IN2(req_out_jump_input_datapath), .Q(and4resu_input_datapath) );

    MUX21X1 U1071(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[36:0][3]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U1072(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[36:0][4]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U1073(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[36:0][5]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U1074(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[36:0][6]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U1075(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[36:0][7]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U1076(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[36:0][8]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U1077(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[36:0][9]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U1078(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[36:0][10]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U1079(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[36:0][11]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U1080(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[36:0][12]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U1081(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[36:0][13]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U1082(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[36:0][14]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U1083(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[36:0][15]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U1084(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[36:0][16]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U1085(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[36:0][17]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U1086(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[36:0][18]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U1087(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[36:0][19]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U1088(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[36:0][20]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U1089(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[36:0][21]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U1090(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[36:0][22]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U1091(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[36:0][23]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U1092(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[36:0][24]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U1093(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[36:0][25]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U1094(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[36:0][26]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U1095(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[36:0][27]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U1096(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[36:0][28]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U1097(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[36:0][29]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U1098(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[36:0][30]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U1099(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[36:0][31]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U1100(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[36:0][32]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U1101(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[36:0][33]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U1102(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[36:0][34]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U1103(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[36:0][35]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U1104(.IN1(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[36:0][36]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U1105(.IN1(int_req_v[36:0][0]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath * 37)]), .S(and4resu_input_datapath), .Q(int_req_v[36:0][0]));
	MUX21X1 U1106(.IN1(int_req_v[36:0][1]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+1]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+1]));
	MUX21X1 U1107(.IN1(int_req_v[36:0][2]),.IN2(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+2]), .S(and4resu_input_datapath), .Q(to_output_req_in_jump_input_datapathput_datapath[(vc_ch_act_out_input_datapath*37)+2]));
	MUX21X1 U1108(.IN1(to_output_resp_input_datapath[vc_ch_act_out_input_datapath]),.IN2(int_resp_v[1:0]), .S(and4resu_input_datapath), .Q(to_output_resp_input_datapath[vc_ch_act_out_input_datapath]));
	MUX21X1 U1109(.IN1(to_output_resp_input_datapath[vc_ch_act_out_input_datapath+1]),.IN2(int_resp_v[1:0]), .S(and4resu_input_datapath), .Q(to_output_resp_input_datapath[vc_ch_act_out_input_datapath+1]));


	BUFX1 U1110 ( .A(read_ptr_ff_fifomodule11[0]), .Y(next_read_ptr_fifomodule11[0]) );
	BUFX1 U1111 ( .A(read_ptr_ff_fifomodule11[1]), .Y(next_read_ptr_fifomodule11[1]) );
	BUFX1 U1112 ( .A(write_ptr_ff_fifomodule11[0]), .Y(next_write_ptr_fifomodule11[0]) );
	BUFX1 U1113 ( .A(write_ptr_ff_fifomodule11[1]), .Y(next_write_ptr_fifomodule11[1]) );

	XNOR2X1 U1114 ( .IN1(write_ptr_ff_fifomodule11[0]), .IN2(read_ptr_ff_fifomodule11[0]), .Q(u1temp_fifomodule11) );
	XNOR2X1 U1115 ( .IN1(write_ptr_ff_fifomodule11[1]), .IN2(read_ptr_ff_fifomodule11[1]), .Q(u2temp_fifomodule11) );
	AND2X1 U1116 ( .A(u1temp_fifomodule11), .B(u2temp_fifomodule11), .Y(empty_vc_buffer11) );
	XOR2X1 U1117 ( .A(write_ptr_ff_fifomodule11[1]), .B(read_ptr_ff_fifomodule11[1]), .Y(u4temp_fifomodule11) );
	AND2X1 U1118 ( .A(u1temp_fifomodule11), .B(u4temp_fifomodule11), .Y(full_vc_buffer11) );
	MUX21X1 U1119 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][0]));
	MUX21X1 U1120 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][1]));
	MUX21X1 U1121 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][2]));
	MUX21X1 U1122 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][3]));
	MUX21X1 U1123 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][4]));
	MUX21X1 U1124 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][5]));
	MUX21X1 U1125 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][6]));
	MUX21X1 U1126 (.IN1(fifo_ff_fifomodule11[read_ptr_ff_fifomodule11[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer11), .Q(to_output_req_in_jump_input_datapath1put_datapath1[36:3][7]));

	INVX1 U1127 ( .A(full_vc_buffer11), .Y(full_vc_buffer11_not_fifomodule) );
	AND2X1 U1128 ( .A(write_flit11_vc_buffer1), .B(full_vc_buffer11_not_fifomodule), .Y(u7temp_fifomodule11) );
	MUX21X1 U1129 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule11), .Q(u9temp_fifomodule11));
	HADDX1 U1130 ( .A0(write_ptr_ff_fifomodule11[0]), .B0(u9temp_fifomodule11), .C1(u10carry_fifomodule11), .SO(next_write_ptr_fifomodule11[0]) );
	HADDX1 U1131 ( .A0(u10carry_fifomodule11), .B0(write_ptr_ff_fifomodule11[1]), .C1(u11carry_fifomodule11), .SO(next_write_ptr_fifomodule11[1]) );

	INVX1 U1132 ( .A(empty_vc_buffer11), .Y(empty_vc_buffer11_not_fifomodule) );
	AND2X1 U1133 ( .A(read_flit11_vc_buffer1), .B(empty_vc_buffer11_not_fifomodule), .Y(u13temp_fifomodule11) );
	MUX21X1 U1134 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule11), .Q(u14temp_fifomodule11));
	HADDX1 U1135 ( .A0(read_ptr_ff_fifomodule11[0]), .B0(u14temp_fifomodule11), .C1(u15carry_fifomodule11), .SO(next_read_ptr_fifomodule11[0]) );
	HADDX1 U1136 ( .A0(u15carry_fifomodule11), .B0(read_ptr_ff_fifomodule11[1]), .C1(u16carry_fifomodule11), .SO(next_read_ptr_fifomodule11[1]) );

	AND2X1 U1137 ( .A(write_flit11_vc_buffer1), .B(full_vc_buffer11), .Y(u17res_fifomodule11) );
	AND2X1 U1138 ( .A(read_flit11_vc_buffer1), .B(empty_vc_buffer11), .Y(u18res_fifomodule11) );
    OR2X1 U1139 ( .A(u17res_fifomodule11), .B(u18res_fifomodule11), .Y(error_vc_buffer11) );
	XOR2X1 U1140 ( .A(write_ptr_ff_fifomodule11[0]), .B(read_ptr_ff_fifomodule11[0]), .Y(fifo_ocup_fifomodule11[0]) );
	INVX1 U1141 ( .A(write_ptr_ff_fifomodule11[0]), .Y(write_ptr_ff_fifomodule11_0_not1) );
	AND2X1 U1142 ( .A(write_ptr_ff_fifomodule11_0_not1), .B(read_ptr_ff_fifomodule11[0]), .Y(b0wire_fifomodule11) );
	XOR2X1 U1143 ( .A(write_ptr_ff_fifomodule11[1]), .B(read_ptr_ff_fifomodule11[1]), .Y(u23temp_fifomodule11) );
	INVX1 U1144 ( .A(write_ptr_ff_fifomodule11[1]), .Y(write_ptr_ff_fifomodule11_1_not1) );
	AND2X1 U1145 ( .A(read_ptr_ff_fifomodule11[1]), .B(write_ptr_ff_fifomodule11_1_not1), .Y(boutb_fifomodule11) );
	XOR2X1 U1146 ( .A(u23temp_fifomodule11), .B(b0wire_fifomodule11), .Y(fifo_ocup_fifomodule11[1]) );
	INVX1 U1147 ( .A(u23temp_fifomodule11), .Y(u23temp_fifomodule11_not_fifomodule11) );
	AND2X1 U1148 ( .A(b0wire_fifomodule11), .B(u23temp_fifomodule11_not_fifomodule11), .Y(bouta_fifomodule11) );
	OR2X1 U1149 ( .A(bouta_fifomodule11), .B(boutb_fifomodule11), .Y(boutmain_fifomodule11) );
	DFFX2 U1150 ( .CLK(clk), .D(fifo_ocup_fifomodule11[0]), .Q(ocup_o[0]) );
	DFFX2 U1151 ( .CLK(clk), .D(fifo_ocup_fifomodule11[1]), .Q(ocup_o[1]) );
	DFFX2 U1152 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule11) );
	DFFX2 U1153 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule11) );
	DFFX2 U1154 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(write_ptr_ff_fifomodule11[0]) );
	DFFX2 U1155 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(read_ptr_ff_fifomodule11[0]) );
	DFFX2 U1156 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(fifo_ff_fifomodule11[0]) );
	DFFX2 U1157 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(write_ptr_ff_fifomodule11[1]) );
	DFFX2 U1158 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(read_ptr_ff_fifomodule11[1]) );
	DFFX2 U1159 ( .CLK(arst_value_fifomodule11), .D(1'b0), .Q(fifo_ff_fifomodule11[1]) );

	DFFX2 U1160 ( .CLK(clk), .D(next_write_ptr_fifomodule11[0]), .Q(write_ptr_ff_fifomodule11[0]) );
	DFFX2 U1161 ( .CLK(clk), .D(next_write_ptr_fifomodule11[1]), .Q(write_ptr_ff_fifomodule11[1]) );
	DFFX2 U1162 ( .CLK(clk), .D(next_read_ptr_fifomodule11[0]), .Q(read_ptr_ff_fifomodule11[0]) );
	DFFX2 U1163 ( .CLK(clk), .D(next_read_ptr_fifomodule11[1]), .Q(read_ptr_ff_fifomodule11[1]) );
	  

	DFFX2 U1164 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][0]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8]) );
	DFFX2 U1165 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][1]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+1]) );
	DFFX2 U1166 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][2]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+2]) );
	DFFX2 U1167 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][3]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+3]) );
	DFFX2 U1168 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][4]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+4]) );
	DFFX2 U1169 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][5]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+5]) );
	DFFX2 U1170 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][6]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+6]) );
	DFFX2 U1171 ( .CLK(u7temp_fifomodule11), .D(from_input_req_in_jump_input_datapath1put_datapath1[36:3][7]), .Q(fifo_ff_fifomodule11[write_ptr_ff_fifomodule11[0]*8+7]) );

    BUFX1 U1172 ( .A(locked_by_route_ff_vc_buffer11), .Y(next_locked_vc_buffer11) );
    BUFX1 U1173(.A(flit11[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][0]));
	BUFX1 U1174(.A(flit11[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][1]));
	BUFX1 U1175(.A(flit11[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][2]));
	BUFX1 U1176(.A(flit11[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][3]));
	BUFX1 U1177(.A(flit11[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][4]));
	BUFX1 U1178(.A(flit11[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][5]));
	BUFX1 U1179(.A(flit11[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][6]));
	BUFX1 U1180(.A(flit11[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][7]));
	BUFX1 U1181(.A(flit11[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][8]));
	BUFX1 U1182(.A(flit11[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][9]));
	BUFX1 U1183(.A(flit11[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][10]));
	BUFX1 U1184(.A(flit11[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][11]));
	BUFX1 U1185(.A(flit11[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][12]));
	BUFX1 U1186(.A(flit11[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][13]));
	BUFX1 U1187(.A(flit11[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][14]));
	BUFX1 U1188(.A(flit11[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][15]));
	BUFX1 U1189(.A(flit11[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][16]));
	BUFX1 U1190(.A(flit11[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][17]));
	BUFX1 U1191(.A(flit11[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][18]));
	BUFX1 U1192(.A(flit11[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][19]));
	BUFX1 U1193(.A(flit11[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][20]));
	BUFX1 U1194(.A(flit11[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][21]));
	BUFX1 U1195(.A(flit11[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][22]));
	BUFX1 U1196(.A(flit11[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][23]));
	BUFX1 U1197(.A(flit11[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][24]));
	BUFX1 U1198(.A(flit11[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][25]));
	BUFX1 U1199(.A(flit11[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][26]));
	BUFX1 U1200(.A(flit11[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][27]));
	BUFX1 U1201(.A(flit11[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][28]));
	BUFX1 U1202(.A(flit11[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][29]));
	BUFX1 U1203(.A(flit11[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][30]));
	BUFX1 U1204(.A(flit11[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][31]));
	BUFX1 U1205(.A(flit11[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][32]));
	BUFX1 U1206(.A(flit11[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[36:3][33]));
    NOR2X1 U1207 ( .IN1(flit11[33]), .IN2(flit11[32]), .QN(norres_vc_buffer11_vc_buffer11) );
    OR4X1 U1208 ( .IN1(flit11[29]), .IN2(flit11[28]), .IN3(flit11[27]), .IN4(flit11[26]), .Y(or1res_vc_buffer11) );
    OR4X1 U1209 ( .IN1(flit11[25]), .IN2(flit11[24]), .IN3(flit11[23]), .IN4(flit11[22]), .Y(or2res_vc_buffer11) );
    OR2X1 U1210 ( .A(or1res_vc_buffer11), .B(or2res_vc_buffer11), .Y(orres_vc_buffer11) );
    AND3X1 U1211 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(norres_vc_buffer11_vc_buffer11), .IN3(orres_vc_buffer11), .Q(finres1_vc_buffer11) );
    MUX21X1 U1212 (.IN1(next_locked_vc_buffer11), .IN2(1'b1), .S(finres1_vc_buffer11), .Q(next_locked_vc_buffer11);
    AND3X1 U1213 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(flit11[33]), .IN3(flit11[32]), .Q(andres1_vc_buffer11) );
    MUX21X1 U1214 (.IN1(next_locked_vc_buffer11), .IN2(1'b0), .S(andres1_vc_buffer11), .Q(next_locked_vc_buffer11);

    INVX1 U1215 ( .A(full_vc_buffer11), .Y(full_vc_buffer11_not) );
    INVX1 U1216 ( .A(locked_by_route_ff_vc_buffer11), .Y(locked_by_route_ff_vc_buffer11_not) );

    MUX21X1 U1217 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer11_not), .S(norres_vc_buffer11_vc_buffer11), .Q(thirdand_vc_buffer11);
    AND3X1 U1218 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[0]), .IN2(full_vc_buffer11_not), .IN3(thirdand_vc_buffer11), .Q(write_flit11_vc_buffer1) );
    AND2X1 U1219 ( .IN1(full_vc_buffer11_not), .IN2(norres_vc_buffer11_vc_buffer11), .Q(from_input_resp_input_datapath1[0]) );
    INVX1 U1220 ( .A(empty_vc_buffer11), .Y(to_output_req_in_jump_input_datapath1put_datapath1[0]) );
    AND2X1 U1221 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[0]), .IN2(to_output_resp_input_datapath1[0]), .Q(read_flit11_vc_buffer1) );
	BUFX1 U1222(.A(to_output_req_in_jump_input_datapath1put_datapath1[2:1]), .Y(2'b00));

	DFFX2 U1223 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1224 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1225 (.IN1(next_locked_vc_buffer11), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer11);

	BUFX1 U1226 ( .A(read_ptr_ff_fifomodule111[0]), .Y(next_read_ptr_fifomodule111[0]) );
	BUFX1 U1227 ( .A(read_ptr_ff_fifomodule111[1]), .Y(next_read_ptr_fifomodule111[1]) );
	BUFX1 U1228 ( .A(write_ptr_ff_fifomodule111[0]), .Y(next_write_ptr_fifomodule111[0]) );
	BUFX1 U1229 ( .A(write_ptr_ff_fifomodule111[1]), .Y(next_write_ptr_fifomodule111[1]) );

	XNOR2X1 U1230 ( .IN1(write_ptr_ff_fifomodule111[0]), .IN2(read_ptr_ff_fifomodule111[0]), .Q(u1temp_fifomodule111) );
	XNOR2X1 U1231 ( .IN1(write_ptr_ff_fifomodule111[1]), .IN2(read_ptr_ff_fifomodule111[1]), .Q(u2temp_fifomodule111) );
	AND2X1 U1232 ( .A(u1temp_fifomodule111), .B(u2temp_fifomodule111), .Y(empty_vc_buffer111) );
	XOR2X1 U1233 ( .A(write_ptr_ff_fifomodule111[1]), .B(read_ptr_ff_fifomodule111[1]), .Y(u4temp_fifomodule111) );
	AND2X1 U1234 ( .A(u1temp_fifomodule111), .B(u4temp_fifomodule111), .Y(full_vc_buffer111) );
	MUX21X1 U1235 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][0]));
	MUX21X1 U1236 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][1]));
	MUX21X1 U1237 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][2]));
	MUX21X1 U1238 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][3]));
	MUX21X1 U1239 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][4]));
	MUX21X1 U1240 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][5]));
	MUX21X1 U1241 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][6]));
	MUX21X1 U1242 (.IN1(fifo_ff_fifomodule111[read_ptr_ff_fifomodule111[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer111), .Q(to_output_req_in_jump_input_datapath1put_datapath1[73:40][7]));

	INVX1 U1243 ( .A(full_vc_buffer111), .Y(full_vc_buffer111_not1_fifomodule1) );
	AND2X1 U1244 ( .A(write_flit111_vc_buffer11), .B(full_vc_buffer111_not1_fifomodule1), .Y(u7temp_fifomodule111) );
	MUX21X1 U1245 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule111), .Q(u9temp_fifomodule111));
	HADDX1 U1246 ( .A0(write_ptr_ff_fifomodule111[0]), .B0(u9temp_fifomodule111), .C1(u10carry_fifomodule111), .SO(next_write_ptr_fifomodule111[0]) );
	HADDX1 U1247 ( .A0(u10carry_fifomodule111), .B0(write_ptr_ff_fifomodule111[1]), .C1(u11carry_fifomodule111), .SO(next_write_ptr_fifomodule111[1]) );

	INVX1 U1248 ( .A(empty_vc_buffer111), .Y(empty_vc_buffer111_not_fifomodule1) );
	AND2X1 U1249 ( .A(read_flit111_vc_buffer11), .B(empty_vc_buffer111_not_fifomodule1), .Y(u13temp_fifomodule111) );
	MUX21X1 U1250 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule111), .Q(u14temp_fifomodule111));
	HADDX1 U1251 ( .A0(read_ptr_ff_fifomodule111[0]), .B0(u14temp_fifomodule111), .C1(u15carry_fifomodule111), .SO(next_read_ptr_fifomodule111[0]) );
	HADDX1 U1252 ( .A0(u15carry_fifomodule111), .B0(read_ptr_ff_fifomodule111[1]), .C1(u16carry_fifomodule111), .SO(next_read_ptr_fifomodule111[1]) );

	AND2X1 U1253 ( .A(write_flit111_vc_buffer11), .B(full_vc_buffer111), .Y(u17res_fifomodule111) );
	AND2X1 U1254 ( .A(read_flit111_vc_buffer11), .B(empty_vc_buffer111), .Y(u18res_fifomodule111) );
    OR2X1 U1255 ( .A(u17res_fifomodule111), .B(u18res_fifomodule111), .Y(error_vc_buffer111) );
	XOR2X1 U1256 ( .A(write_ptr_ff_fifomodule111[0]), .B(read_ptr_ff_fifomodule111[0]), .Y(fifo_ocup_fifomodule111[0]) );
	INVX1 U1257 ( .A(write_ptr_ff_fifomodule111[0]), .Y(write_ptr_ff_fifomodule111_0_not11) );
	AND2X1 U1258 ( .A(write_ptr_ff_fifomodule111_0_not11), .B(read_ptr_ff_fifomodule111[0]), .Y(b0wire_fifomodule111) );
	XOR2X1 U1259 ( .A(write_ptr_ff_fifomodule111[1]), .B(read_ptr_ff_fifomodule111[1]), .Y(u23temp_fifomodule111) );
	INVX1 U1260 ( .A(write_ptr_ff_fifomodule111[1]), .Y(write_ptr_ff_fifomodule111_1_not11) );
	AND2X1 U1261 ( .A(read_ptr_ff_fifomodule111[1]), .B(write_ptr_ff_fifomodule111_1_not11), .Y(boutb_fifomodule111) );
	XOR2X1 U1262 ( .A(u23temp_fifomodule111), .B(b0wire_fifomodule111), .Y(fifo_ocup_fifomodule111[1]) );
	INVX1 U1263 ( .A(u23temp_fifomodule111), .Y(u23temp_fifomodule111_not_fifomodule1) );
	AND2X1 U1264 ( .A(b0wire_fifomodule111), .B(u23temp_fifomodule111_not_fifomodule1), .Y(bouta_fifomodule111) );
	OR2X1 U1265 ( .A(bouta_fifomodule111), .B(boutb_fifomodule111), .Y(boutmain_fifomodule111) );
	DFFX2 U1266 ( .CLK(clk), .D(fifo_ocup_fifomodule111[0]), .Q(ocup_o[0]) );
	DFFX2 U1267 ( .CLK(clk), .D(fifo_ocup_fifomodule111[1]), .Q(ocup_o[1]) );
	DFFX2 U1268 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule111) );
	DFFX2 U1269 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule111) );
	DFFX2 U1270 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(write_ptr_ff_fifomodule111[0]) );
	DFFX2 U1271 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(read_ptr_ff_fifomodule111[0]) );
	DFFX2 U1272 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(fifo_ff_fifomodule111[0]) );
	DFFX2 U1273 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(write_ptr_ff_fifomodule111[1]) );
	DFFX2 U1274 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(read_ptr_ff_fifomodule111[1]) );
	DFFX2 U1275 ( .CLK(arst_value_fifomodule111), .D(1'b0), .Q(fifo_ff_fifomodule111[1]) );

	DFFX2 U1276 ( .CLK(clk), .D(next_write_ptr_fifomodule111[0]), .Q(write_ptr_ff_fifomodule111[0]) );
	DFFX2 U1277 ( .CLK(clk), .D(next_write_ptr_fifomodule111[1]), .Q(write_ptr_ff_fifomodule111[1]) );
	DFFX2 U1278 ( .CLK(clk), .D(next_read_ptr_fifomodule111[0]), .Q(read_ptr_ff_fifomodule111[0]) );
	DFFX2 U1279 ( .CLK(clk), .D(next_read_ptr_fifomodule111[1]), .Q(read_ptr_ff_fifomodule111[1]) );
	  

	DFFX2 U1280 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][0]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8]) );
	DFFX2 U1281 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][1]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+1]) );
	DFFX2 U1282 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][2]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+2]) );
	DFFX2 U1283 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][3]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+3]) );
	DFFX2 U1284 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][4]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+4]) );
	DFFX2 U1285 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][5]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+5]) );
	DFFX2 U1286 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][6]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+6]) );
	DFFX2 U1287 ( .CLK(u7temp_fifomodule111), .D(from_input_req_in_jump_input_datapath1put_datapath1[73:40][7]), .Q(fifo_ff_fifomodule111[write_ptr_ff_fifomodule111[0]*8+7]) );

    BUFX1 U1288 ( .A(locked_by_route_ff_vc_buffer111), .Y(next_locked_vc_buffer111) );
    BUFX1 U1289(.A(flit111[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][0]));
	BUFX1 U1290(.A(flit111[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][1]));
	BUFX1 U1291(.A(flit111[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][2]));
	BUFX1 U1292(.A(flit111[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][3]));
	BUFX1 U1293(.A(flit111[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][4]));
	BUFX1 U1294(.A(flit111[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][5]));
	BUFX1 U1295(.A(flit111[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][6]));
	BUFX1 U1296(.A(flit111[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][7]));
	BUFX1 U1297(.A(flit111[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][8]));
	BUFX1 U1298(.A(flit111[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][9]));
	BUFX1 U1299(.A(flit111[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][10]));
	BUFX1 U1300(.A(flit111[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][11]));
	BUFX1 U1301(.A(flit111[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][12]));
	BUFX1 U1302(.A(flit111[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][13]));
	BUFX1 U1303(.A(flit111[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][14]));
	BUFX1 U1304(.A(flit111[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][15]));
	BUFX1 U1305(.A(flit111[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][16]));
	BUFX1 U1306(.A(flit111[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][17]));
	BUFX1 U1307(.A(flit111[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][18]));
	BUFX1 U1308(.A(flit111[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][19]));
	BUFX1 U1309(.A(flit111[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][20]));
	BUFX1 U1310(.A(flit111[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][21]));
	BUFX1 U1311(.A(flit111[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][22]));
	BUFX1 U1312(.A(flit111[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][23]));
	BUFX1 U1313(.A(flit111[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][24]));
	BUFX1 U1314(.A(flit111[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][25]));
	BUFX1 U1315(.A(flit111[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][26]));
	BUFX1 U1316(.A(flit111[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][27]));
	BUFX1 U1317(.A(flit111[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][28]));
	BUFX1 U1318(.A(flit111[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][29]));
	BUFX1 U1319(.A(flit111[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][30]));
	BUFX1 U1320(.A(flit111[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][31]));
	BUFX1 U1321(.A(flit111[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][32]));
	BUFX1 U1322(.A(flit111[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[73:40][33]));
    NOR2X1 U1323 ( .IN1(flit111[33]), .IN2(flit111[32]), .QN(norres_vc_buffer111_vc_buffer1) );
    OR4X1 U1324 ( .IN1(flit111[29]), .IN2(flit111[28]), .IN3(flit111[27]), .IN4(flit111[26]), .Y(or1res_vc_buffer111) );
    OR4X1 U1325 ( .IN1(flit111[25]), .IN2(flit111[24]), .IN3(flit111[23]), .IN4(flit111[22]), .Y(or2res_vc_buffer111) );
    OR2X1 U1326 ( .A(or1res_vc_buffer111), .B(or2res_vc_buffer111), .Y(orres_vc_buffer111) );
    AND3X1 U1327 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(norres_vc_buffer111_vc_buffer1), .IN3(orres_vc_buffer111), .Q(finres1_vc_buffer111) );
    MUX21X1 U1328 (.IN1(next_locked_vc_buffer111), .IN2(1'b1), .S(finres1_vc_buffer111), .Q(next_locked_vc_buffer111);
    AND3X1 U1329 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(flit111[33]), .IN3(flit111[32]), .Q(andres1_vc_buffer111) );
    MUX21X1 U1330 (.IN1(next_locked_vc_buffer111), .IN2(1'b0), .S(andres1_vc_buffer111), .Q(next_locked_vc_buffer111);

    INVX1 U1331 ( .A(full_vc_buffer111), .Y(full_vc_buffer111_not1) );
    INVX1 U1332 ( .A(locked_by_route_ff_vc_buffer111), .Y(locked_by_route_ff_vc_buffer111_not1) );

    MUX21X1 U1333 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer111_not1), .S(norres_vc_buffer111_vc_buffer1), .Q(thirdand_vc_buffer111);
    AND3X1 U1334 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[37]), .IN2(full_vc_buffer111_not1), .IN3(thirdand_vc_buffer111), .Q(write_flit111_vc_buffer11) );
    AND2X1 U1335 ( .IN1(full_vc_buffer111_not1), .IN2(norres_vc_buffer111_vc_buffer1), .Q(from_input_resp_input_datapath1[1]) );
    INVX1 U1336 ( .A(empty_vc_buffer111), .Y(to_output_req_in_jump_input_datapath1put_datapath1[37]) );
    AND2X1 U1337 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[37]), .IN2(to_output_resp_input_datapath1[1]), .Q(read_flit111_vc_buffer11) );
	BUFX1 U1338(.A(to_output_req_in_jump_input_datapath1put_datapath1[39:38]), .Y(2'b01));

	DFFX2 U1339 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1340 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1341 (.IN1(next_locked_vc_buffer111), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer111);


	BUFX1 U1342 ( .A(read_ptr_ff_fifomodule112[0]), .Y(next_read_ptr_fifomodule112[0]) );
	BUFX1 U1343 ( .A(read_ptr_ff_fifomodule112[1]), .Y(next_read_ptr_fifomodule112[1]) );
	BUFX1 U1344 ( .A(write_ptr_ff_fifomodule112[0]), .Y(next_write_ptr_fifomodule112[0]) );
	BUFX1 U1345 ( .A(write_ptr_ff_fifomodule112[1]), .Y(next_write_ptr_fifomodule112[1]) );

	XNOR2X1 U1346 ( .IN1(write_ptr_ff_fifomodule112[0]), .IN2(read_ptr_ff_fifomodule112[0]), .Q(u1temp_fifomodule112) );
	XNOR2X1 U1347 ( .IN1(write_ptr_ff_fifomodule112[1]), .IN2(read_ptr_ff_fifomodule112[1]), .Q(u2temp_fifomodule112) );
	AND2X1 U1348 ( .A(u1temp_fifomodule112), .B(u2temp_fifomodule112), .Y(empty_vc_buffer112) );
	XOR2X1 U1349 ( .A(write_ptr_ff_fifomodule112[1]), .B(read_ptr_ff_fifomodule112[1]), .Y(u4temp_fifomodule112) );
	AND2X1 U1350 ( .A(u1temp_fifomodule112), .B(u4temp_fifomodule112), .Y(full_vc_buffer112) );
	MUX21X1 U1351 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][0]));
	MUX21X1 U1352 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][1]));
	MUX21X1 U1353 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][2]));
	MUX21X1 U1354 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][3]));
	MUX21X1 U1355 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][4]));
	MUX21X1 U1356 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][5]));
	MUX21X1 U1357 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][6]));
	MUX21X1 U1358 (.IN1(fifo_ff_fifomodule112[read_ptr_ff_fifomodule112[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer112), .Q(to_output_req_in_jump_input_datapath1put_datapath1[110:77][7]));

	INVX1 U1359 ( .A(full_vc_buffer112), .Y(full_vc_buffer112_not2_fifomodule2) );
	AND2X1 U1360 ( .A(write_flit112_vc_buffer21), .B(full_vc_buffer112_not2_fifomodule2), .Y(u7temp_fifomodule112) );
	MUX21X1 U1361 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule112), .Q(u9temp_fifomodule112));
	HADDX1 U1362 ( .A0(write_ptr_ff_fifomodule112[0]), .B0(u9temp_fifomodule112), .C1(u10carry_fifomodule112), .SO(next_write_ptr_fifomodule112[0]) );
	HADDX1 U1363 ( .A0(u10carry_fifomodule112), .B0(write_ptr_ff_fifomodule112[1]), .C1(u11carry_fifomodule112), .SO(next_write_ptr_fifomodule112[1]) );

	INVX1 U1364 ( .A(empty_vc_buffer112), .Y(empty_vc_buffer112_not_fifomodule2) );
	AND2X1 U1365 ( .A(read_flit112_vc_buffer21), .B(empty_vc_buffer112_not_fifomodule2), .Y(u13temp_fifomodule112) );
	MUX21X1 U1366 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule112), .Q(u14temp_fifomodule112));
	HADDX1 U1367 ( .A0(read_ptr_ff_fifomodule112[0]), .B0(u14temp_fifomodule112), .C1(u15carry_fifomodule112), .SO(next_read_ptr_fifomodule112[0]) );
	HADDX1 U1368 ( .A0(u15carry_fifomodule112), .B0(read_ptr_ff_fifomodule112[1]), .C1(u16carry_fifomodule112), .SO(next_read_ptr_fifomodule112[1]) );

	AND2X1 U1369 ( .A(write_flit112_vc_buffer21), .B(full_vc_buffer112), .Y(u17res_fifomodule112) );
	AND2X1 U1370 ( .A(read_flit112_vc_buffer21), .B(empty_vc_buffer112), .Y(u18res_fifomodule112) );
    OR2X1 U1371 ( .A(u17res_fifomodule112), .B(u18res_fifomodule112), .Y(error_vc_buffer112) );
	XOR2X1 U1372 ( .A(write_ptr_ff_fifomodule112[0]), .B(read_ptr_ff_fifomodule112[0]), .Y(fifo_ocup_fifomodule112[0]) );
	INVX1 U1373 ( .A(write_ptr_ff_fifomodule112[0]), .Y(write_ptr_ff_fifomodule112_0_not21) );
	AND2X1 U1374 ( .A(write_ptr_ff_fifomodule112_0_not21), .B(read_ptr_ff_fifomodule112[0]), .Y(b0wire_fifomodule112) );
	XOR2X1 U1375 ( .A(write_ptr_ff_fifomodule112[1]), .B(read_ptr_ff_fifomodule112[1]), .Y(u23temp_fifomodule112) );
	INVX1 U1376 ( .A(write_ptr_ff_fifomodule112[1]), .Y(write_ptr_ff_fifomodule112_1_not21) );
	AND2X1 U1377 ( .A(read_ptr_ff_fifomodule112[1]), .B(write_ptr_ff_fifomodule112_1_not21), .Y(boutb_fifomodule112) );
	XOR2X1 U1378 ( .A(u23temp_fifomodule112), .B(b0wire_fifomodule112), .Y(fifo_ocup_fifomodule112[1]) );
	INVX1 U1379 ( .A(u23temp_fifomodule112), .Y(u23temp_fifomodule112_not_fifomodule2) );
	AND2X1 U1380 ( .A(b0wire_fifomodule112), .B(u23temp_fifomodule112_not_fifomodule2), .Y(bouta_fifomodule112) );
	OR2X1 U1381 ( .A(bouta_fifomodule112), .B(boutb_fifomodule112), .Y(boutmain_fifomodule112) );
	DFFX2 U1382 ( .CLK(clk), .D(fifo_ocup_fifomodule112[0]), .Q(ocup_o[0]) );
	DFFX2 U1383 ( .CLK(clk), .D(fifo_ocup_fifomodule112[1]), .Q(ocup_o[1]) );
	DFFX2 U1384 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule112) );
	DFFX2 U1385 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule112) );
	DFFX2 U1386 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(write_ptr_ff_fifomodule112[0]) );
	DFFX2 U1387 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(read_ptr_ff_fifomodule112[0]) );
	DFFX2 U1388 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(fifo_ff_fifomodule112[0]) );
	DFFX2 U1389 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(write_ptr_ff_fifomodule112[1]) );
	DFFX2 U1390 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(read_ptr_ff_fifomodule112[1]) );
	DFFX2 U1391 ( .CLK(arst_value_fifomodule112), .D(1'b0), .Q(fifo_ff_fifomodule112[1]) );

	DFFX2 U1392 ( .CLK(clk), .D(next_write_ptr_fifomodule112[0]), .Q(write_ptr_ff_fifomodule112[0]) );
	DFFX2 U1393 ( .CLK(clk), .D(next_write_ptr_fifomodule112[1]), .Q(write_ptr_ff_fifomodule112[1]) );
	DFFX2 U1394 ( .CLK(clk), .D(next_read_ptr_fifomodule112[0]), .Q(read_ptr_ff_fifomodule112[0]) );
	DFFX2 U1395 ( .CLK(clk), .D(next_read_ptr_fifomodule112[1]), .Q(read_ptr_ff_fifomodule112[1]) );
	  

	DFFX2 U1396 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][0]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8]) );
	DFFX2 U1397 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][1]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+1]) );
	DFFX2 U1398 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][2]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+2]) );
	DFFX2 U1399 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][3]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+3]) );
	DFFX2 U1400 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][4]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+4]) );
	DFFX2 U1401 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][5]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+5]) );
	DFFX2 U1402 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][6]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+6]) );
	DFFX2 U1403 ( .CLK(u7temp_fifomodule112), .D(from_input_req_in_jump_input_datapath1put_datapath1[110:77][7]), .Q(fifo_ff_fifomodule112[write_ptr_ff_fifomodule112[0]*8+7]) );

    BUFX1 U1404 ( .A(locked_by_route_ff_vc_buffer112), .Y(next_locked_vc_buffer112) );
    BUFX1 U1405(.A(flit112[0]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][0]));
	BUFX1 U1406(.A(flit112[1]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][1]));
	BUFX1 U1407(.A(flit112[2]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][2]));
	BUFX1 U1408(.A(flit112[3]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][3]));
	BUFX1 U1409(.A(flit112[4]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][4]));
	BUFX1 U1410(.A(flit112[5]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][5]));
	BUFX1 U1411(.A(flit112[6]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][6]));
	BUFX1 U1412(.A(flit112[7]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][7]));
	BUFX1 U1413(.A(flit112[8]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][8]));
	BUFX1 U1414(.A(flit112[9]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][9]));
	BUFX1 U1415(.A(flit112[10]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][10]));
	BUFX1 U1416(.A(flit112[11]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][11]));
	BUFX1 U1417(.A(flit112[12]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][12]));
	BUFX1 U1418(.A(flit112[13]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][13]));
	BUFX1 U1419(.A(flit112[14]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][14]));
	BUFX1 U1420(.A(flit112[15]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][15]));
	BUFX1 U1421(.A(flit112[16]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][16]));
	BUFX1 U1422(.A(flit112[17]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][17]));
	BUFX1 U1423(.A(flit112[18]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][18]));
	BUFX1 U1424(.A(flit112[19]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][19]));
	BUFX1 U1425(.A(flit112[20]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][20]));
	BUFX1 U1426(.A(flit112[21]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][21]));
	BUFX1 U1427(.A(flit112[22]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][22]));
	BUFX1 U1428(.A(flit112[23]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][23]));
	BUFX1 U1429(.A(flit112[24]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][24]));
	BUFX1 U1430(.A(flit112[25]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][25]));
	BUFX1 U1431(.A(flit112[26]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][26]));
	BUFX1 U1432(.A(flit112[27]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][27]));
	BUFX1 U1433(.A(flit112[28]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][28]));
	BUFX1 U1434(.A(flit112[29]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][29]));
	BUFX1 U1435(.A(flit112[30]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][30]));
	BUFX1 U1436(.A(flit112[31]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][31]));
	BUFX1 U1437(.A(flit112[32]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][32]));
	BUFX1 U1438(.A(flit112[33]), .Y(from_input_req_in_jump_input_datapath1put_datapath1[110:77][33]));
    NOR2X1 U1439 ( .IN1(flit112[33]), .IN2(flit112[32]), .QN(norres_vc_buffer112_vc_buffer2) );
    OR4X1 U1440 ( .IN1(flit112[29]), .IN2(flit112[28]), .IN3(flit112[27]), .IN4(flit112[26]), .Y(or1res_vc_buffer112) );
    OR4X1 U1441 ( .IN1(flit112[25]), .IN2(flit112[24]), .IN3(flit112[23]), .IN4(flit112[22]), .Y(or2res_vc_buffer112) );
    OR2X1 U1442 ( .A(or1res_vc_buffer112), .B(or2res_vc_buffer112), .Y(orres_vc_buffer112) );
    AND3X1 U1443 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(norres_vc_buffer112_vc_buffer2), .IN3(orres_vc_buffer112), .Q(finres1_vc_buffer112) );
    MUX21X1 U1444 (.IN1(next_locked_vc_buffer112), .IN2(1'b1), .S(finres1_vc_buffer112), .Q(next_locked_vc_buffer112);
    AND3X1 U1445 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(flit112[33]), .IN3(flit112[32]), .Q(andres1_vc_buffer112) );
    MUX21X1 U1446 (.IN1(next_locked_vc_buffer112), .IN2(1'b0), .S(andres1_vc_buffer112), .Q(next_locked_vc_buffer112);

    INVX1 U1447 ( .A(full_vc_buffer112), .Y(full_vc_buffer112_not2) );
    INVX1 U1448 ( .A(locked_by_route_ff_vc_buffer112), .Y(locked_by_route_ff_vc_buffer112_not2) );

    MUX21X1 U1449 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer112_not2), .S(norres_vc_buffer112_vc_buffer2), .Q(thirdand_vc_buffer112);
    AND3X1 U1450 ( .IN1(from_input_req_in_jump_input_datapath1put_datapath1[74]), .IN2(full_vc_buffer112_not2), .IN3(thirdand_vc_buffer112), .Q(write_flit112_vc_buffer21) );
    AND2X1 U1451 ( .IN1(full_vc_buffer112_not2), .IN2(norres_vc_buffer112_vc_buffer2), .Q(from_input_resp_input_datapath1[2]) );
    INVX1 U1452 ( .A(empty_vc_buffer112), .Y(to_output_req_in_jump_input_datapath1put_datapath1[74]) );
    AND2X1 U1453 ( .IN1(to_output_req_in_jump_input_datapath1put_datapath1[74]), .IN2(to_output_resp_input_datapath1[2]), .Q(read_flit112_vc_buffer21) );
	BUFX1 U1454(.A(to_output_req_in_jump_input_datapath1put_datapath1[76:75]), .Y(2'b10));

	DFFX2 U1455 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1456 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1457 (.IN1(next_locked_vc_buffer112), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer112);

	BUFX1 U1458(.A(from_input_req_in_jump_input_datapath1put_datapath1[77]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U1459(.A(from_input_req_in_jump_input_datapath1put_datapath1[78]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U1460(.A(from_input_req_in_jump_input_datapath1put_datapath1[79]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U1461(.A(from_input_req_in_jump_input_datapath1put_datapath1[80]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U1462(.A(from_input_req_in_jump_input_datapath1put_datapath1[81]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U1463(.A(from_input_req_in_jump_input_datapath1put_datapath1[82]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U1464(.A(from_input_req_in_jump_input_datapath1put_datapath1[83]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U1465(.A(from_input_req_in_jump_input_datapath1put_datapath1[84]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U1466(.A(from_input_req_in_jump_input_datapath1put_datapath1[85]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U1467(.A(from_input_req_in_jump_input_datapath1put_datapath1[86]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U1468(.A(from_input_req_in_jump_input_datapath1put_datapath1[87]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U1469(.A(from_input_req_in_jump_input_datapath1put_datapath1[88]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U1470(.A(from_input_req_in_jump_input_datapath1put_datapath1[89]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U1471(.A(from_input_req_in_jump_input_datapath1put_datapath1[90]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U1472(.A(from_input_req_in_jump_input_datapath1put_datapath1[91]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U1473(.A(from_input_req_in_jump_input_datapath1put_datapath1[92]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U1474(.A(from_input_req_in_jump_input_datapath1put_datapath1[93]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U1475(.A(from_input_req_in_jump_input_datapath1put_datapath1[94]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U1476(.A(from_input_req_in_jump_input_datapath1put_datapath1[95]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U1477(.A(from_input_req_in_jump_input_datapath1put_datapath1[96]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U1478(.A(from_input_req_in_jump_input_datapath1put_datapath1[97]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U1479(.A(from_input_req_in_jump_input_datapath1put_datapath1[98]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U1480(.A(from_input_req_in_jump_input_datapath1put_datapath1[99]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U1481(.A(from_input_req_in_jump_input_datapath1put_datapath1[100]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U1482(.A(from_input_req_in_jump_input_datapath1put_datapath1[101]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U1483(.A(from_input_req_in_jump_input_datapath1put_datapath1[102]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U1484(.A(from_input_req_in_jump_input_datapath1put_datapath1[103]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U1485(.A(from_input_req_in_jump_input_datapath1put_datapath1[104]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U1486(.A(from_input_req_in_jump_input_datapath1put_datapath1[105]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U1487(.A(from_input_req_in_jump_input_datapath1put_datapath1[106]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U1488(.A(from_input_req_in_jump_input_datapath1put_datapath1[107]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U1489(.A(from_input_req_in_jump_input_datapath1put_datapath1[108]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U1490(.A(from_input_req_in_jump_input_datapath1put_datapath1[109]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U1491(.A(from_input_req_in_jump_input_datapath1put_datapath1[110]), .Y(ext_req_v_i[73:37][36]));
    XNOR2X1 U1492 ( .IN1(ext_req_v_i[73:37][1]), .IN2(i_input_datapath1[0]), .QN(xnor1resu_input_datapath1) );
    XNOR2X1 U1493 ( .IN1(ext_req_v_i[73:37][2]), .IN2(i_input_datapath1[1]), .QN(xnor2resu_input_datapath1) );
    AND2X1 U1494 ( .IN1(xnor1resu_input_datapath1), .IN2(xnor2resu_input_datapath1), .Q(and1resu_input_datapath1) );
    AND3X1 U1495 ( .IN1(and1resu_input_datapath1), .IN2(ext_req_v_i[73:37][0]), .IN2(ext_req_v_i[73:37][0]), .Q(cond1line_input_datapath1) );
    MUX21X1 U1496 (.IN1(vc_ch_act_in_input_datapath1[0]), .IN2(i_input_datapath1[0]), .S(cond1line_input_datapath1), .Q(vc_ch_act_in_input_datapath1[0]));
    MUX21X1 U1497 (.IN1(vc_ch_act_in_input_datapath1[1]), .IN2(i_input_datapath1[1]), .S(cond1line_input_datapath1), .Q(vc_ch_act_in_input_datapath1[1]));
    MUX21X1 U1498 (.IN1(req_in_jump_input_datapath1), .IN2(1), .S(cond1line_input_datapath1), .Q(req_in_jump_input_datapath1));
	BUFX1 U1499(.A(from_input_req_in_jump_input_datapath1put_datapath1[40]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U1500(.A(from_input_req_in_jump_input_datapath1put_datapath1[41]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U1501(.A(from_input_req_in_jump_input_datapath1put_datapath1[42]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U1502(.A(from_input_req_in_jump_input_datapath1put_datapath1[43]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U1503(.A(from_input_req_in_jump_input_datapath1put_datapath1[44]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U1504(.A(from_input_req_in_jump_input_datapath1put_datapath1[45]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U1505(.A(from_input_req_in_jump_input_datapath1put_datapath1[46]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U1506(.A(from_input_req_in_jump_input_datapath1put_datapath1[47]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U1507(.A(from_input_req_in_jump_input_datapath1put_datapath1[48]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U1508(.A(from_input_req_in_jump_input_datapath1put_datapath1[49]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U1509(.A(from_input_req_in_jump_input_datapath1put_datapath1[50]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U1510(.A(from_input_req_in_jump_input_datapath1put_datapath1[51]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U1511(.A(from_input_req_in_jump_input_datapath1put_datapath1[52]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U1512(.A(from_input_req_in_jump_input_datapath1put_datapath1[53]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U1513(.A(from_input_req_in_jump_input_datapath1put_datapath1[54]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U1514(.A(from_input_req_in_jump_input_datapath1put_datapath1[55]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U1515(.A(from_input_req_in_jump_input_datapath1put_datapath1[56]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U1516(.A(from_input_req_in_jump_input_datapath1put_datapath1[57]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U1517(.A(from_input_req_in_jump_input_datapath1put_datapath1[58]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U1518(.A(from_input_req_in_jump_input_datapath1put_datapath1[59]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U1519(.A(from_input_req_in_jump_input_datapath1put_datapath1[60]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U1520(.A(from_input_req_in_jump_input_datapath1put_datapath1[61]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U1521(.A(from_input_req_in_jump_input_datapath1put_datapath1[62]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U1522(.A(from_input_req_in_jump_input_datapath1put_datapath1[63]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U1523(.A(from_input_req_in_jump_input_datapath1put_datapath1[64]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U1524(.A(from_input_req_in_jump_input_datapath1put_datapath1[65]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U1525(.A(from_input_req_in_jump_input_datapath1put_datapath1[66]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U1526(.A(from_input_req_in_jump_input_datapath1put_datapath1[67]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U1527(.A(from_input_req_in_jump_input_datapath1put_datapath1[68]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U1528(.A(from_input_req_in_jump_input_datapath1put_datapath1[69]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U1529(.A(from_input_req_in_jump_input_datapath1put_datapath1[70]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U1530(.A(from_input_req_in_jump_input_datapath1put_datapath1[71]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U1531(.A(from_input_req_in_jump_input_datapath1put_datapath1[72]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U1532(.A(from_input_req_in_jump_input_datapath1put_datapath1[73]), .Y(ext_req_v_i[73:37][36]));

	BUFX1 U1533(.A(from_input_req_in_jump_input_datapath1put_datapath1[3]), .Y(ext_req_v_i[73:37][3]));
	BUFX1 U1534(.A(from_input_req_in_jump_input_datapath1put_datapath1[4]), .Y(ext_req_v_i[73:37][4]));
	BUFX1 U1535(.A(from_input_req_in_jump_input_datapath1put_datapath1[5]), .Y(ext_req_v_i[73:37][5]));
	BUFX1 U1536(.A(from_input_req_in_jump_input_datapath1put_datapath1[6]), .Y(ext_req_v_i[73:37][6]));
	BUFX1 U1537(.A(from_input_req_in_jump_input_datapath1put_datapath1[7]), .Y(ext_req_v_i[73:37][7]));
	BUFX1 U1538(.A(from_input_req_in_jump_input_datapath1put_datapath1[8]), .Y(ext_req_v_i[73:37][8]));
	BUFX1 U1539(.A(from_input_req_in_jump_input_datapath1put_datapath1[9]), .Y(ext_req_v_i[73:37][9]));
	BUFX1 U1540(.A(from_input_req_in_jump_input_datapath1put_datapath1[10]), .Y(ext_req_v_i[73:37][10]));
	BUFX1 U1541(.A(from_input_req_in_jump_input_datapath1put_datapath1[11]), .Y(ext_req_v_i[73:37][11]));
	BUFX1 U1542(.A(from_input_req_in_jump_input_datapath1put_datapath1[12]), .Y(ext_req_v_i[73:37][12]));
	BUFX1 U1543(.A(from_input_req_in_jump_input_datapath1put_datapath1[13]), .Y(ext_req_v_i[73:37][13]));
	BUFX1 U1544(.A(from_input_req_in_jump_input_datapath1put_datapath1[14]), .Y(ext_req_v_i[73:37][14]));
	BUFX1 U1545(.A(from_input_req_in_jump_input_datapath1put_datapath1[15]), .Y(ext_req_v_i[73:37][15]));
	BUFX1 U1546(.A(from_input_req_in_jump_input_datapath1put_datapath1[16]), .Y(ext_req_v_i[73:37][16]));
	BUFX1 U1547(.A(from_input_req_in_jump_input_datapath1put_datapath1[17]), .Y(ext_req_v_i[73:37][17]));
	BUFX1 U1548(.A(from_input_req_in_jump_input_datapath1put_datapath1[18]), .Y(ext_req_v_i[73:37][18]));
	BUFX1 U1549(.A(from_input_req_in_jump_input_datapath1put_datapath1[19]), .Y(ext_req_v_i[73:37][19]));
	BUFX1 U1550(.A(from_input_req_in_jump_input_datapath1put_datapath1[20]), .Y(ext_req_v_i[73:37][20]));
	BUFX1 U1551(.A(from_input_req_in_jump_input_datapath1put_datapath1[21]), .Y(ext_req_v_i[73:37][21]));
	BUFX1 U1552(.A(from_input_req_in_jump_input_datapath1put_datapath1[22]), .Y(ext_req_v_i[73:37][22]));
	BUFX1 U1553(.A(from_input_req_in_jump_input_datapath1put_datapath1[23]), .Y(ext_req_v_i[73:37][23]));
	BUFX1 U1554(.A(from_input_req_in_jump_input_datapath1put_datapath1[24]), .Y(ext_req_v_i[73:37][24]));
	BUFX1 U1555(.A(from_input_req_in_jump_input_datapath1put_datapath1[25]), .Y(ext_req_v_i[73:37][25]));
	BUFX1 U1556(.A(from_input_req_in_jump_input_datapath1put_datapath1[26]), .Y(ext_req_v_i[73:37][26]));
	BUFX1 U1557(.A(from_input_req_in_jump_input_datapath1put_datapath1[27]), .Y(ext_req_v_i[73:37][27]));
	BUFX1 U1558(.A(from_input_req_in_jump_input_datapath1put_datapath1[28]), .Y(ext_req_v_i[73:37][28]));
	BUFX1 U1559(.A(from_input_req_in_jump_input_datapath1put_datapath1[29]), .Y(ext_req_v_i[73:37][29]));
	BUFX1 U1560(.A(from_input_req_in_jump_input_datapath1put_datapath1[30]), .Y(ext_req_v_i[73:37][30]));
	BUFX1 U1561(.A(from_input_req_in_jump_input_datapath1put_datapath1[31]), .Y(ext_req_v_i[73:37][31]));
	BUFX1 U1562(.A(from_input_req_in_jump_input_datapath1put_datapath1[32]), .Y(ext_req_v_i[73:37][32]));
	BUFX1 U1563(.A(from_input_req_in_jump_input_datapath1put_datapath1[33]), .Y(ext_req_v_i[73:37][33]));
	BUFX1 U1564(.A(from_input_req_in_jump_input_datapath1put_datapath1[34]), .Y(ext_req_v_i[73:37][34]));
	BUFX1 U1565(.A(from_input_req_in_jump_input_datapath1put_datapath1[35]), .Y(ext_req_v_i[73:37][35]));
	BUFX1 U1566(.A(from_input_req_in_jump_input_datapath1put_datapath1[36]), .Y(ext_req_v_i[73:37][36]));

    MUX21X1 U1567 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1 * 37]), .IN2(ext_req_v_i[73:37][0]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1 * 37]));
    MUX21X1 U1568 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+2]), .IN2(vc_ch_act_in_input_datapath1[1]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+2]));
    MUX21X1 U1569 (.IN1(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+1]), .IN2(vc_ch_act_in_input_datapath1[0]), .S(req_in_jump_input_datapath1), .Q(from_input_req_in_jump_input_datapath1put_datapath1[vc_ch_act_in_input_datapath1*37+1]));
    MUX21X1 U1570 (.IN1(ext_resp_v_o[2:1][0]), .IN2(from_input_resp_input_datapath1[vc_ch_act_in_input_datapath1]), .S(req_in_jump_input_datapath1), .Q(ext_resp_v_o[2:1][0]));

    INVX1 U1571 ( .A(req_in_jump_input_datapath1), .Y(req_in_jump_input_datapath1_not) );
    MUX21X1 U1572 (.IN1(ext_resp_v_o[2:1][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath1_not), .Q(ext_resp_v_o[2:1][0]));
    BUFX1 U1573(.A(from_input_req_in_jump_input_datapath1put_datapath1[34]), .Y(ext_req_v_i[73:37][34]));

    XOR2X1 U1574 ( .IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b1), .Q(xor1resu_input_datapath1) );
    MUX21X1 U1575 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(xor1resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U1576 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b0), .S(xor1resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[1]));
    AND2X1 U1577 ( .IN1(xor1resu_input_datapath1), .IN2(to_output_req_in_jump_input_datapath1put_datapath1[j_input_datapath1*37]), .Q(and2resu_input_datapath1) );
    MUX21X1 U1578 (.IN1(vc_ch_act_out_input_datapath1[0]), .IN2(j_input_datapath1[0]), .S(and2resu_input_datapath1), .Q(vc_ch_act_out_input_datapath1[0]));
    MUX21X1 U1579 (.IN1(vc_ch_act_out_input_datapath1[1]), .IN2(j_input_datapath1[1]), .S(and2resu_input_datapath1), .Q(vc_ch_act_out_input_datapath1[1]));
    MUX21X1 U1580 (.IN1(req_out_jump_input_datapath1), .IN2(1'b1), .S(and2resu_input_datapath1), .Q(req_out_jump_input_datapath1));
    MUX21X1 U1581 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(and2resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U1582 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b1), .S(and2resu_input_datapath1), .Q(_sv2v_jump_input_datapath1[1]));
    HADDX1 U1583 ( .A0(j_input_datapath1[0]), .B0(1'b1), .C1(j_input_datapath1[1]), .SO(j_input_datapath1[0]) );
    HADDX1 U1584 ( .A0(j_input_datapath1[0]), .B0(1'b1), .C1(j_input_datapath1[1]), .SO(j_input_datapath1[0]) );
    AND2X1 U1585 ( .IN1(xor1resu_input_datapath1), .IN2(to_output_req_in_jump_input_datapath1put_datapath1[j_input_datapath1*37]), .Q(and3resu) );
    NAND2X1 U1586(.A(_sv2v_jump_input_datapath1[0]),.B(_sv2v_jump_input_datapath1[1]),.Y(nand1resu_input_datapath11));
    MUX21X1 U1587 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(1'b0), .S(nand1resu_input_datapath11), .Q(_sv2v_jump_input_datapath1[0]));
    MUX21X1 U1588 (.IN1(_sv2v_jump_input_datapath1[1]), .IN2(1'b0), .S(nand1resu_input_datapath11), .Q(_sv2v_jump_input_datapath1[1]));
    XNOR2X1 U1589 (.IN1(_sv2v_jump_input_datapath1[0]), .IN2(_sv2v_jump_input_datapath1[1]), .Q(xnor23resu_input_datapath1) );
    AND2X1 U1590 ( .IN1(xnor23resu_input_datapath1), .IN2(req_out_jump_input_datapath1), .Q(and4resu_input_datapath1) );

    MUX21X1 U1591(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[73:37][3]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U1592(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[73:37][4]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U1593(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[73:37][5]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U1594(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[73:37][6]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U1595(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[73:37][7]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U1596(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[73:37][8]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U1597(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[73:37][9]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U1598(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[73:37][10]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U1599(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[73:37][11]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U1600(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[73:37][12]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U1601(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[73:37][13]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U1602(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[73:37][14]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U1603(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[73:37][15]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U1604(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[73:37][16]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U1605(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[73:37][17]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U1606(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[73:37][18]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U1607(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[73:37][19]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U1608(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[73:37][20]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U1609(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[73:37][21]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U1610(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[73:37][22]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U1611(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[73:37][23]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U1612(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[73:37][24]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U1613(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[73:37][25]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U1614(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[73:37][26]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U1615(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[73:37][27]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U1616(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[73:37][28]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U1617(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[73:37][29]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U1618(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[73:37][30]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U1619(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[73:37][31]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U1620(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[73:37][32]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U1621(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[73:37][33]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U1622(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[73:37][34]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U1623(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[73:37][35]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U1624(.IN1(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[73:37][36]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U1625(.IN1(int_req_v[73:37][0]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1 * 37)]), .S(and4resu_input_datapath1), .Q(int_req_v[73:37][0]));
	MUX21X1 U1626(.IN1(int_req_v[73:37][1]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+1]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+1]));
	MUX21X1 U1627(.IN1(int_req_v[73:37][2]),.IN2(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+2]), .S(and4resu_input_datapath1), .Q(to_output_req_in_jump_input_datapath1put_datapath1[(vc_ch_act_out_input_datapath1*37)+2]));
	MUX21X1 U1628(.IN1(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1]),.IN2(int_resp_v[2:1]), .S(and4resu_input_datapath1), .Q(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1]));
	MUX21X1 U1629(.IN1(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1+1]),.IN2(int_resp_v[2:1]), .S(and4resu_input_datapath1), .Q(to_output_resp_input_datapath1[vc_ch_act_out_input_datapath1+1]));

	BUFX1 U1630 ( .A(read_ptr_ff_fifomodule22[0]), .Y(next_read_ptr_fifomodule22[0]) );
	BUFX1 U1631 ( .A(read_ptr_ff_fifomodule22[1]), .Y(next_read_ptr_fifomodule22[1]) );
	BUFX1 U1632 ( .A(write_ptr_ff_fifomodule22[0]), .Y(next_write_ptr_fifomodule22[0]) );
	BUFX1 U1633 ( .A(write_ptr_ff_fifomodule22[1]), .Y(next_write_ptr_fifomodule22[1]) );

	XNOR2X1 U1634 ( .IN1(write_ptr_ff_fifomodule22[0]), .IN2(read_ptr_ff_fifomodule22[0]), .Q(u1temp_fifomodule22) );
	XNOR2X1 U1635 ( .IN1(write_ptr_ff_fifomodule22[1]), .IN2(read_ptr_ff_fifomodule22[1]), .Q(u2temp_fifomodule22) );
	AND2X1 U1636 ( .A(u1temp_fifomodule22), .B(u2temp_fifomodule22), .Y(empty_vc_buffer22) );
	XOR2X1 U1637 ( .A(write_ptr_ff_fifomodule22[1]), .B(read_ptr_ff_fifomodule22[1]), .Y(u4temp_fifomodule22) );
	AND2X1 U1638 ( .A(u1temp_fifomodule22), .B(u4temp_fifomodule22), .Y(full_vc_buffer22) );
	MUX21X1 U1639 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][0]));
	MUX21X1 U1640 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][1]));
	MUX21X1 U1641 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][2]));
	MUX21X1 U1642 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][3]));
	MUX21X1 U1643 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][4]));
	MUX21X1 U1644 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][5]));
	MUX21X1 U1645 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][6]));
	MUX21X1 U1646 (.IN1(fifo_ff_fifomodule22[read_ptr_ff_fifomodule22[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer22), .Q(to_output_req_in_jump_input_datapath2put_datapath2[36:3][7]));

	INVX1 U1647 ( .A(full_vc_buffer22), .Y(full_vc_buffer22_not_fifomodule) );
	AND2X1 U1648 ( .A(write_flit22_vc_buffer2), .B(full_vc_buffer22_not_fifomodule), .Y(u7temp_fifomodule22) );
	MUX21X1 U1649 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule22), .Q(u9temp_fifomodule22));
	HADDX1 U1650 ( .A0(write_ptr_ff_fifomodule22[0]), .B0(u9temp_fifomodule22), .C1(u10carry_fifomodule22), .SO(next_write_ptr_fifomodule22[0]) );
	HADDX1 U1651 ( .A0(u10carry_fifomodule22), .B0(write_ptr_ff_fifomodule22[1]), .C1(u11carry_fifomodule22), .SO(next_write_ptr_fifomodule22[1]) );

	INVX1 U1652 ( .A(empty_vc_buffer22), .Y(empty_vc_buffer22_not_fifomodule) );
	AND2X1 U1653 ( .A(read_flit22_vc_buffer2), .B(empty_vc_buffer22_not_fifomodule), .Y(u13temp_fifomodule22) );
	MUX21X1 U1654 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule22), .Q(u14temp_fifomodule22));
	HADDX1 U1655 ( .A0(read_ptr_ff_fifomodule22[0]), .B0(u14temp_fifomodule22), .C1(u15carry_fifomodule22), .SO(next_read_ptr_fifomodule22[0]) );
	HADDX1 U1656 ( .A0(u15carry_fifomodule22), .B0(read_ptr_ff_fifomodule22[1]), .C1(u16carry_fifomodule22), .SO(next_read_ptr_fifomodule22[1]) );

	AND2X1 U1657 ( .A(write_flit22_vc_buffer2), .B(full_vc_buffer22), .Y(u17res_fifomodule22) );
	AND2X1 U1658 ( .A(read_flit22_vc_buffer2), .B(empty_vc_buffer22), .Y(u18res_fifomodule22) );
    OR2X1 U1659 ( .A(u17res_fifomodule22), .B(u18res_fifomodule22), .Y(error_vc_buffer22) );
	XOR2X1 U1660 ( .A(write_ptr_ff_fifomodule22[0]), .B(read_ptr_ff_fifomodule22[0]), .Y(fifo_ocup_fifomodule22[0]) );
	INVX1 U1661 ( .A(write_ptr_ff_fifomodule22[0]), .Y(write_ptr_ff_fifomodule22_0_not2) );
	AND2X1 U1662 ( .A(write_ptr_ff_fifomodule22_0_not2), .B(read_ptr_ff_fifomodule22[0]), .Y(b0wire_fifomodule22) );
	XOR2X1 U1663 ( .A(write_ptr_ff_fifomodule22[1]), .B(read_ptr_ff_fifomodule22[1]), .Y(u23temp_fifomodule22) );
	INVX1 U1664 ( .A(write_ptr_ff_fifomodule22[1]), .Y(write_ptr_ff_fifomodule22_1_not2) );
	AND2X1 U1665 ( .A(read_ptr_ff_fifomodule22[1]), .B(write_ptr_ff_fifomodule22_1_not2), .Y(boutb_fifomodule22) );
	XOR2X1 U1666 ( .A(u23temp_fifomodule22), .B(b0wire_fifomodule22), .Y(fifo_ocup_fifomodule22[1]) );
	INVX1 U1667 ( .A(u23temp_fifomodule22), .Y(u23temp_fifomodule22_not_fifomodule22) );
	AND2X1 U1668 ( .A(b0wire_fifomodule22), .B(u23temp_fifomodule22_not_fifomodule22), .Y(bouta_fifomodule22) );
	OR2X1 U1669 ( .A(bouta_fifomodule22), .B(boutb_fifomodule22), .Y(boutmain_fifomodule22) );
	DFFX2 U1670 ( .CLK(clk), .D(fifo_ocup_fifomodule22[0]), .Q(ocup_o[0]) );
	DFFX2 U1671 ( .CLK(clk), .D(fifo_ocup_fifomodule22[1]), .Q(ocup_o[1]) );
	DFFX2 U1672 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule22) );
	DFFX2 U1673 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule22) );
	DFFX2 U1674 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(write_ptr_ff_fifomodule22[0]) );
	DFFX2 U1675 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(read_ptr_ff_fifomodule22[0]) );
	DFFX2 U1676 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(fifo_ff_fifomodule22[0]) );
	DFFX2 U1677 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(write_ptr_ff_fifomodule22[1]) );
	DFFX2 U1678 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(read_ptr_ff_fifomodule22[1]) );
	DFFX2 U1679 ( .CLK(arst_value_fifomodule22), .D(1'b0), .Q(fifo_ff_fifomodule22[1]) );

	DFFX2 U1680 ( .CLK(clk), .D(next_write_ptr_fifomodule22[0]), .Q(write_ptr_ff_fifomodule22[0]) );
	DFFX2 U1681 ( .CLK(clk), .D(next_write_ptr_fifomodule22[1]), .Q(write_ptr_ff_fifomodule22[1]) );
	DFFX2 U1682 ( .CLK(clk), .D(next_read_ptr_fifomodule22[0]), .Q(read_ptr_ff_fifomodule22[0]) );
	DFFX2 U1683 ( .CLK(clk), .D(next_read_ptr_fifomodule22[1]), .Q(read_ptr_ff_fifomodule22[1]) );
	  

	DFFX2 U1684 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][0]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8]) );
	DFFX2 U1685 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][1]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+1]) );
	DFFX2 U1686 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][2]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+2]) );
	DFFX2 U1687 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][3]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+3]) );
	DFFX2 U1688 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][4]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+4]) );
	DFFX2 U1689 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][5]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+5]) );
	DFFX2 U1690 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][6]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+6]) );
	DFFX2 U1691 ( .CLK(u7temp_fifomodule22), .D(from_input_req_in_jump_input_datapath2put_datapath2[36:3][7]), .Q(fifo_ff_fifomodule22[write_ptr_ff_fifomodule22[0]*8+7]) );

    BUFX1 U1692 ( .A(locked_by_route_ff_vc_buffer22), .Y(next_locked_vc_buffer22) );
    BUFX1 U1693(.A(flit22[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][0]));
	BUFX1 U1694(.A(flit22[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][1]));
	BUFX1 U1695(.A(flit22[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][2]));
	BUFX1 U1696(.A(flit22[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][3]));
	BUFX1 U1697(.A(flit22[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][4]));
	BUFX1 U1698(.A(flit22[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][5]));
	BUFX1 U1699(.A(flit22[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][6]));
	BUFX1 U1700(.A(flit22[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][7]));
	BUFX1 U1701(.A(flit22[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][8]));
	BUFX1 U1702(.A(flit22[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][9]));
	BUFX1 U1703(.A(flit22[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][10]));
	BUFX1 U1704(.A(flit22[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][11]));
	BUFX1 U1705(.A(flit22[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][12]));
	BUFX1 U1706(.A(flit22[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][13]));
	BUFX1 U1707(.A(flit22[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][14]));
	BUFX1 U1708(.A(flit22[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][15]));
	BUFX1 U1709(.A(flit22[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][16]));
	BUFX1 U1710(.A(flit22[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][17]));
	BUFX1 U1711(.A(flit22[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][18]));
	BUFX1 U1712(.A(flit22[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][19]));
	BUFX1 U1713(.A(flit22[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][20]));
	BUFX1 U1714(.A(flit22[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][21]));
	BUFX1 U1715(.A(flit22[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][22]));
	BUFX1 U1716(.A(flit22[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][23]));
	BUFX1 U1717(.A(flit22[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][24]));
	BUFX1 U1718(.A(flit22[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][25]));
	BUFX1 U1719(.A(flit22[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][26]));
	BUFX1 U1720(.A(flit22[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][27]));
	BUFX1 U1721(.A(flit22[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][28]));
	BUFX1 U1722(.A(flit22[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][29]));
	BUFX1 U1723(.A(flit22[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][30]));
	BUFX1 U1724(.A(flit22[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][31]));
	BUFX1 U1725(.A(flit22[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][32]));
	BUFX1 U1726(.A(flit22[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[36:3][33]));
    NOR2X1 U1727 ( .IN1(flit22[33]), .IN2(flit22[32]), .QN(norres_vc_buffer22_vc_buffer22) );
    OR4X1 U1728 ( .IN1(flit22[29]), .IN2(flit22[28]), .IN3(flit22[27]), .IN4(flit22[26]), .Y(or1res_vc_buffer22) );
    OR4X1 U1729 ( .IN1(flit22[25]), .IN2(flit22[24]), .IN3(flit22[23]), .IN4(flit22[22]), .Y(or2res_vc_buffer22) );
    OR2X1 U1730 ( .A(or1res_vc_buffer22), .B(or2res_vc_buffer22), .Y(orres_vc_buffer22) );
    AND3X1 U1731 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(norres_vc_buffer22_vc_buffer22), .IN3(orres_vc_buffer22), .Q(finres1_vc_buffer22) );
    MUX21X1 U1732 (.IN1(next_locked_vc_buffer22), .IN2(1'b1), .S(finres1_vc_buffer22), .Q(next_locked_vc_buffer22);
    AND3X1 U1733 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(flit22[33]), .IN3(flit22[32]), .Q(andres1_vc_buffer22) );
    MUX21X1 U1734 (.IN1(next_locked_vc_buffer22), .IN2(1'b0), .S(andres1_vc_buffer22), .Q(next_locked_vc_buffer22);

    INVX1 U1735 ( .A(full_vc_buffer22), .Y(full_vc_buffer22_not) );
    INVX1 U1736 ( .A(locked_by_route_ff_vc_buffer22), .Y(locked_by_route_ff_vc_buffer22_not) );

    MUX21X1 U1737 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer22_not), .S(norres_vc_buffer22_vc_buffer22), .Q(thirdand_vc_buffer22);
    AND3X1 U1738 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[0]), .IN2(full_vc_buffer22_not), .IN3(thirdand_vc_buffer22), .Q(write_flit22_vc_buffer2) );
    AND2X1 U1739 ( .IN1(full_vc_buffer22_not), .IN2(norres_vc_buffer22_vc_buffer22), .Q(from_input_resp_input_datapath2[0]) );
    INVX1 U1740 ( .A(empty_vc_buffer22), .Y(to_output_req_in_jump_input_datapath2put_datapath2[0]) );
    AND2X1 U1741 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[0]), .IN2(to_output_resp_input_datapath2[0]), .Q(read_flit22_vc_buffer2) );
	BUFX1 U1742(.A(to_output_req_in_jump_input_datapath2put_datapath2[2:1]), .Y(2'b00));

	DFFX2 U1743 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1744 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1745 (.IN1(next_locked_vc_buffer22), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer22);

	BUFX1 U1746 ( .A(read_ptr_ff_fifomodule221[0]), .Y(next_read_ptr_fifomodule221[0]) );
	BUFX1 U1747 ( .A(read_ptr_ff_fifomodule221[1]), .Y(next_read_ptr_fifomodule221[1]) );
	BUFX1 U1748 ( .A(write_ptr_ff_fifomodule221[0]), .Y(next_write_ptr_fifomodule221[0]) );
	BUFX1 U1749 ( .A(write_ptr_ff_fifomodule221[1]), .Y(next_write_ptr_fifomodule221[1]) );

	XNOR2X1 U1750 ( .IN1(write_ptr_ff_fifomodule221[0]), .IN2(read_ptr_ff_fifomodule221[0]), .Q(u1temp_fifomodule221) );
	XNOR2X1 U1751 ( .IN1(write_ptr_ff_fifomodule221[1]), .IN2(read_ptr_ff_fifomodule221[1]), .Q(u2temp_fifomodule221) );
	AND2X1 U1752 ( .A(u1temp_fifomodule221), .B(u2temp_fifomodule221), .Y(empty_vc_buffer221) );
	XOR2X1 U1753 ( .A(write_ptr_ff_fifomodule221[1]), .B(read_ptr_ff_fifomodule221[1]), .Y(u4temp_fifomodule221) );
	AND2X1 U1754 ( .A(u1temp_fifomodule221), .B(u4temp_fifomodule221), .Y(full_vc_buffer221) );
	MUX21X1 U1755 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][0]));
	MUX21X1 U1756 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][1]));
	MUX21X1 U1757 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][2]));
	MUX21X1 U1758 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][3]));
	MUX21X1 U1759 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][4]));
	MUX21X1 U1760 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][5]));
	MUX21X1 U1761 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][6]));
	MUX21X1 U1762 (.IN1(fifo_ff_fifomodule221[read_ptr_ff_fifomodule221[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer221), .Q(to_output_req_in_jump_input_datapath2put_datapath2[73:40][7]));

	INVX1 U1763 ( .A(full_vc_buffer221), .Y(full_vc_buffer221_not1_fifomodule1) );
	AND2X1 U1764 ( .A(write_flit221_vc_buffer12), .B(full_vc_buffer221_not1_fifomodule1), .Y(u7temp_fifomodule221) );
	MUX21X1 U1765 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule221), .Q(u9temp_fifomodule221));
	HADDX1 U1766 ( .A0(write_ptr_ff_fifomodule221[0]), .B0(u9temp_fifomodule221), .C1(u10carry_fifomodule221), .SO(next_write_ptr_fifomodule221[0]) );
	HADDX1 U1767 ( .A0(u10carry_fifomodule221), .B0(write_ptr_ff_fifomodule221[1]), .C1(u11carry_fifomodule221), .SO(next_write_ptr_fifomodule221[1]) );

	INVX1 U1768 ( .A(empty_vc_buffer221), .Y(empty_vc_buffer221_not_fifomodule1) );
	AND2X1 U1769 ( .A(read_flit221_vc_buffer12), .B(empty_vc_buffer221_not_fifomodule1), .Y(u13temp_fifomodule221) );
	MUX21X1 U1770 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule221), .Q(u14temp_fifomodule221));
	HADDX1 U1771 ( .A0(read_ptr_ff_fifomodule221[0]), .B0(u14temp_fifomodule221), .C1(u15carry_fifomodule221), .SO(next_read_ptr_fifomodule221[0]) );
	HADDX1 U1772 ( .A0(u15carry_fifomodule221), .B0(read_ptr_ff_fifomodule221[1]), .C1(u16carry_fifomodule221), .SO(next_read_ptr_fifomodule221[1]) );

	AND2X1 U1773 ( .A(write_flit221_vc_buffer12), .B(full_vc_buffer221), .Y(u17res_fifomodule221) );
	AND2X1 U1774 ( .A(read_flit221_vc_buffer12), .B(empty_vc_buffer221), .Y(u18res_fifomodule221) );
    OR2X1 U1775 ( .A(u17res_fifomodule221), .B(u18res_fifomodule221), .Y(error_vc_buffer221) );
	XOR2X1 U1776 ( .A(write_ptr_ff_fifomodule221[0]), .B(read_ptr_ff_fifomodule221[0]), .Y(fifo_ocup_fifomodule221[0]) );
	INVX1 U1777 ( .A(write_ptr_ff_fifomodule221[0]), .Y(write_ptr_ff_fifomodule221_0_not12) );
	AND2X1 U1778 ( .A(write_ptr_ff_fifomodule221_0_not12), .B(read_ptr_ff_fifomodule221[0]), .Y(b0wire_fifomodule221) );
	XOR2X1 U1779 ( .A(write_ptr_ff_fifomodule221[1]), .B(read_ptr_ff_fifomodule221[1]), .Y(u23temp_fifomodule221) );
	INVX1 U1780 ( .A(write_ptr_ff_fifomodule221[1]), .Y(write_ptr_ff_fifomodule221_1_not12) );
	AND2X1 U1781 ( .A(read_ptr_ff_fifomodule221[1]), .B(write_ptr_ff_fifomodule221_1_not12), .Y(boutb_fifomodule221) );
	XOR2X1 U1782 ( .A(u23temp_fifomodule221), .B(b0wire_fifomodule221), .Y(fifo_ocup_fifomodule221[1]) );
	INVX1 U1783 ( .A(u23temp_fifomodule221), .Y(u23temp_fifomodule221_not_fifomodule1) );
	AND2X1 U1784 ( .A(b0wire_fifomodule221), .B(u23temp_fifomodule221_not_fifomodule1), .Y(bouta_fifomodule221) );
	OR2X1 U1785 ( .A(bouta_fifomodule221), .B(boutb_fifomodule221), .Y(boutmain_fifomodule221) );
	DFFX2 U1786 ( .CLK(clk), .D(fifo_ocup_fifomodule221[0]), .Q(ocup_o[0]) );
	DFFX2 U1787 ( .CLK(clk), .D(fifo_ocup_fifomodule221[1]), .Q(ocup_o[1]) );
	DFFX2 U1788 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule221) );
	DFFX2 U1789 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule221) );
	DFFX2 U1790 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(write_ptr_ff_fifomodule221[0]) );
	DFFX2 U1791 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(read_ptr_ff_fifomodule221[0]) );
	DFFX2 U1792 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(fifo_ff_fifomodule221[0]) );
	DFFX2 U1793 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(write_ptr_ff_fifomodule221[1]) );
	DFFX2 U1794 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(read_ptr_ff_fifomodule221[1]) );
	DFFX2 U1795 ( .CLK(arst_value_fifomodule221), .D(1'b0), .Q(fifo_ff_fifomodule221[1]) );

	DFFX2 U1796 ( .CLK(clk), .D(next_write_ptr_fifomodule221[0]), .Q(write_ptr_ff_fifomodule221[0]) );
	DFFX2 U1797 ( .CLK(clk), .D(next_write_ptr_fifomodule221[1]), .Q(write_ptr_ff_fifomodule221[1]) );
	DFFX2 U1798 ( .CLK(clk), .D(next_read_ptr_fifomodule221[0]), .Q(read_ptr_ff_fifomodule221[0]) );
	DFFX2 U1799 ( .CLK(clk), .D(next_read_ptr_fifomodule221[1]), .Q(read_ptr_ff_fifomodule221[1]) );
	  

	DFFX2 U1800 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][0]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8]) );
	DFFX2 U1801 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][1]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+1]) );
	DFFX2 U1802 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][2]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+2]) );
	DFFX2 U1803 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][3]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+3]) );
	DFFX2 U1804 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][4]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+4]) );
	DFFX2 U1805 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][5]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+5]) );
	DFFX2 U1806 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][6]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+6]) );
	DFFX2 U1807 ( .CLK(u7temp_fifomodule221), .D(from_input_req_in_jump_input_datapath2put_datapath2[73:40][7]), .Q(fifo_ff_fifomodule221[write_ptr_ff_fifomodule221[0]*8+7]) );

    BUFX1 U1808 ( .A(locked_by_route_ff_vc_buffer221), .Y(next_locked_vc_buffer221) );
    BUFX1 U1809(.A(flit221[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][0]));
	BUFX1 U1810(.A(flit221[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][1]));
	BUFX1 U1811(.A(flit221[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][2]));
	BUFX1 U1812(.A(flit221[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][3]));
	BUFX1 U1813(.A(flit221[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][4]));
	BUFX1 U1814(.A(flit221[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][5]));
	BUFX1 U1815(.A(flit221[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][6]));
	BUFX1 U1816(.A(flit221[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][7]));
	BUFX1 U1817(.A(flit221[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][8]));
	BUFX1 U1818(.A(flit221[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][9]));
	BUFX1 U1819(.A(flit221[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][10]));
	BUFX1 U1820(.A(flit221[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][11]));
	BUFX1 U1821(.A(flit221[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][12]));
	BUFX1 U1822(.A(flit221[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][13]));
	BUFX1 U1823(.A(flit221[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][14]));
	BUFX1 U1824(.A(flit221[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][15]));
	BUFX1 U1825(.A(flit221[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][16]));
	BUFX1 U1826(.A(flit221[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][17]));
	BUFX1 U1827(.A(flit221[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][18]));
	BUFX1 U1828(.A(flit221[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][19]));
	BUFX1 U1829(.A(flit221[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][20]));
	BUFX1 U1830(.A(flit221[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][21]));
	BUFX1 U1831(.A(flit221[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][22]));
	BUFX1 U1832(.A(flit221[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][23]));
	BUFX1 U1833(.A(flit221[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][24]));
	BUFX1 U1834(.A(flit221[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][25]));
	BUFX1 U1835(.A(flit221[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][26]));
	BUFX1 U1836(.A(flit221[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][27]));
	BUFX1 U1837(.A(flit221[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][28]));
	BUFX1 U1838(.A(flit221[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][29]));
	BUFX1 U1839(.A(flit221[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][30]));
	BUFX1 U1840(.A(flit221[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][31]));
	BUFX1 U1841(.A(flit221[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][32]));
	BUFX1 U1842(.A(flit221[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[73:40][33]));
    NOR2X1 U1843 ( .IN1(flit221[33]), .IN2(flit221[32]), .QN(norres_vc_buffer221_vc_buffer1) );
    OR4X1 U1844 ( .IN1(flit221[29]), .IN2(flit221[28]), .IN3(flit221[27]), .IN4(flit221[26]), .Y(or1res_vc_buffer221) );
    OR4X1 U1845 ( .IN1(flit221[25]), .IN2(flit221[24]), .IN3(flit221[23]), .IN4(flit221[22]), .Y(or2res_vc_buffer221) );
    OR2X1 U1846 ( .A(or1res_vc_buffer221), .B(or2res_vc_buffer221), .Y(orres_vc_buffer221) );
    AND3X1 U1847 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(norres_vc_buffer221_vc_buffer1), .IN3(orres_vc_buffer221), .Q(finres1_vc_buffer221) );
    MUX21X1 U1848 (.IN1(next_locked_vc_buffer221), .IN2(1'b1), .S(finres1_vc_buffer221), .Q(next_locked_vc_buffer221);
    AND3X1 U1849 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(flit221[33]), .IN3(flit221[32]), .Q(andres1_vc_buffer221) );
    MUX21X1 U1850 (.IN1(next_locked_vc_buffer221), .IN2(1'b0), .S(andres1_vc_buffer221), .Q(next_locked_vc_buffer221);

    INVX1 U1851 ( .A(full_vc_buffer221), .Y(full_vc_buffer221_not1) );
    INVX1 U1852 ( .A(locked_by_route_ff_vc_buffer221), .Y(locked_by_route_ff_vc_buffer221_not1) );

    MUX21X1 U1853 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer221_not1), .S(norres_vc_buffer221_vc_buffer1), .Q(thirdand_vc_buffer221);
    AND3X1 U1854 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[37]), .IN2(full_vc_buffer221_not1), .IN3(thirdand_vc_buffer221), .Q(write_flit221_vc_buffer12) );
    AND2X1 U1855 ( .IN1(full_vc_buffer221_not1), .IN2(norres_vc_buffer221_vc_buffer1), .Q(from_input_resp_input_datapath2[1]) );
    INVX1 U1856 ( .A(empty_vc_buffer221), .Y(to_output_req_in_jump_input_datapath2put_datapath2[37]) );
    AND2X1 U1857 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[37]), .IN2(to_output_resp_input_datapath2[1]), .Q(read_flit221_vc_buffer12) );
	BUFX1 U1858(.A(to_output_req_in_jump_input_datapath2put_datapath2[39:38]), .Y(2'b01));

	DFFX2 U1859 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1860 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1861 (.IN1(next_locked_vc_buffer221), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer221);


	BUFX1 U1862 ( .A(read_ptr_ff_fifomodule222[0]), .Y(next_read_ptr_fifomodule222[0]) );
	BUFX1 U1863 ( .A(read_ptr_ff_fifomodule222[1]), .Y(next_read_ptr_fifomodule222[1]) );
	BUFX1 U1864 ( .A(write_ptr_ff_fifomodule222[0]), .Y(next_write_ptr_fifomodule222[0]) );
	BUFX1 U1865 ( .A(write_ptr_ff_fifomodule222[1]), .Y(next_write_ptr_fifomodule222[1]) );

	XNOR2X1 U1866 ( .IN1(write_ptr_ff_fifomodule222[0]), .IN2(read_ptr_ff_fifomodule222[0]), .Q(u1temp_fifomodule222) );
	XNOR2X1 U1867 ( .IN1(write_ptr_ff_fifomodule222[1]), .IN2(read_ptr_ff_fifomodule222[1]), .Q(u2temp_fifomodule222) );
	AND2X1 U1868 ( .A(u1temp_fifomodule222), .B(u2temp_fifomodule222), .Y(empty_vc_buffer222) );
	XOR2X1 U1869 ( .A(write_ptr_ff_fifomodule222[1]), .B(read_ptr_ff_fifomodule222[1]), .Y(u4temp_fifomodule222) );
	AND2X1 U1870 ( .A(u1temp_fifomodule222), .B(u4temp_fifomodule222), .Y(full_vc_buffer222) );
	MUX21X1 U1871 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][0]));
	MUX21X1 U1872 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][1]));
	MUX21X1 U1873 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][2]));
	MUX21X1 U1874 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][3]));
	MUX21X1 U1875 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][4]));
	MUX21X1 U1876 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][5]));
	MUX21X1 U1877 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][6]));
	MUX21X1 U1878 (.IN1(fifo_ff_fifomodule222[read_ptr_ff_fifomodule222[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer222), .Q(to_output_req_in_jump_input_datapath2put_datapath2[110:77][7]));

	INVX1 U1879 ( .A(full_vc_buffer222), .Y(full_vc_buffer222_not2_fifomodule2) );
	AND2X1 U1880 ( .A(write_flit222_vc_buffer22), .B(full_vc_buffer222_not2_fifomodule2), .Y(u7temp_fifomodule222) );
	MUX21X1 U1881 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule222), .Q(u9temp_fifomodule222));
	HADDX1 U1882 ( .A0(write_ptr_ff_fifomodule222[0]), .B0(u9temp_fifomodule222), .C1(u10carry_fifomodule222), .SO(next_write_ptr_fifomodule222[0]) );
	HADDX1 U1883 ( .A0(u10carry_fifomodule222), .B0(write_ptr_ff_fifomodule222[1]), .C1(u11carry_fifomodule222), .SO(next_write_ptr_fifomodule222[1]) );

	INVX1 U1884 ( .A(empty_vc_buffer222), .Y(empty_vc_buffer222_not_fifomodule2) );
	AND2X1 U1885 ( .A(read_flit222_vc_buffer22), .B(empty_vc_buffer222_not_fifomodule2), .Y(u13temp_fifomodule222) );
	MUX21X1 U1886 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule222), .Q(u14temp_fifomodule222));
	HADDX1 U1887 ( .A0(read_ptr_ff_fifomodule222[0]), .B0(u14temp_fifomodule222), .C1(u15carry_fifomodule222), .SO(next_read_ptr_fifomodule222[0]) );
	HADDX1 U1888 ( .A0(u15carry_fifomodule222), .B0(read_ptr_ff_fifomodule222[1]), .C1(u16carry_fifomodule222), .SO(next_read_ptr_fifomodule222[1]) );

	AND2X1 U1889 ( .A(write_flit222_vc_buffer22), .B(full_vc_buffer222), .Y(u17res_fifomodule222) );
	AND2X1 U1890 ( .A(read_flit222_vc_buffer22), .B(empty_vc_buffer222), .Y(u18res_fifomodule222) );
    OR2X1 U1891 ( .A(u17res_fifomodule222), .B(u18res_fifomodule222), .Y(error_vc_buffer222) );
	XOR2X1 U1892 ( .A(write_ptr_ff_fifomodule222[0]), .B(read_ptr_ff_fifomodule222[0]), .Y(fifo_ocup_fifomodule222[0]) );
	INVX1 U1893 ( .A(write_ptr_ff_fifomodule222[0]), .Y(write_ptr_ff_fifomodule222_0_not22) );
	AND2X1 U1894 ( .A(write_ptr_ff_fifomodule222_0_not22), .B(read_ptr_ff_fifomodule222[0]), .Y(b0wire_fifomodule222) );
	XOR2X1 U1895 ( .A(write_ptr_ff_fifomodule222[1]), .B(read_ptr_ff_fifomodule222[1]), .Y(u23temp_fifomodule222) );
	INVX1 U1896 ( .A(write_ptr_ff_fifomodule222[1]), .Y(write_ptr_ff_fifomodule222_1_not22) );
	AND2X1 U1897 ( .A(read_ptr_ff_fifomodule222[1]), .B(write_ptr_ff_fifomodule222_1_not22), .Y(boutb_fifomodule222) );
	XOR2X1 U1898 ( .A(u23temp_fifomodule222), .B(b0wire_fifomodule222), .Y(fifo_ocup_fifomodule222[1]) );
	INVX1 U1899 ( .A(u23temp_fifomodule222), .Y(u23temp_fifomodule222_not_fifomodule2) );
	AND2X1 U1900 ( .A(b0wire_fifomodule222), .B(u23temp_fifomodule222_not_fifomodule2), .Y(bouta_fifomodule222) );
	OR2X1 U1901 ( .A(bouta_fifomodule222), .B(boutb_fifomodule222), .Y(boutmain_fifomodule222) );
	DFFX2 U1902 ( .CLK(clk), .D(fifo_ocup_fifomodule222[0]), .Q(ocup_o[0]) );
	DFFX2 U1903 ( .CLK(clk), .D(fifo_ocup_fifomodule222[1]), .Q(ocup_o[1]) );
	DFFX2 U1904 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule222) );
	DFFX2 U1905 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule222) );
	DFFX2 U1906 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(write_ptr_ff_fifomodule222[0]) );
	DFFX2 U1907 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(read_ptr_ff_fifomodule222[0]) );
	DFFX2 U1908 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(fifo_ff_fifomodule222[0]) );
	DFFX2 U1909 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(write_ptr_ff_fifomodule222[1]) );
	DFFX2 U1910 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(read_ptr_ff_fifomodule222[1]) );
	DFFX2 U1911 ( .CLK(arst_value_fifomodule222), .D(1'b0), .Q(fifo_ff_fifomodule222[1]) );

	DFFX2 U1912 ( .CLK(clk), .D(next_write_ptr_fifomodule222[0]), .Q(write_ptr_ff_fifomodule222[0]) );
	DFFX2 U1913 ( .CLK(clk), .D(next_write_ptr_fifomodule222[1]), .Q(write_ptr_ff_fifomodule222[1]) );
	DFFX2 U1914 ( .CLK(clk), .D(next_read_ptr_fifomodule222[0]), .Q(read_ptr_ff_fifomodule222[0]) );
	DFFX2 U1915 ( .CLK(clk), .D(next_read_ptr_fifomodule222[1]), .Q(read_ptr_ff_fifomodule222[1]) );
	  

	DFFX2 U1916 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][0]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8]) );
	DFFX2 U1917 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][1]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+1]) );
	DFFX2 U1918 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][2]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+2]) );
	DFFX2 U1919 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][3]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+3]) );
	DFFX2 U1920 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][4]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+4]) );
	DFFX2 U1921 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][5]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+5]) );
	DFFX2 U1922 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][6]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+6]) );
	DFFX2 U1923 ( .CLK(u7temp_fifomodule222), .D(from_input_req_in_jump_input_datapath2put_datapath2[110:77][7]), .Q(fifo_ff_fifomodule222[write_ptr_ff_fifomodule222[0]*8+7]) );

    BUFX1 U1924 ( .A(locked_by_route_ff_vc_buffer222), .Y(next_locked_vc_buffer222) );
    BUFX1 U1925(.A(flit222[0]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][0]));
	BUFX1 U1926(.A(flit222[1]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][1]));
	BUFX1 U1927(.A(flit222[2]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][2]));
	BUFX1 U1928(.A(flit222[3]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][3]));
	BUFX1 U1929(.A(flit222[4]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][4]));
	BUFX1 U1930(.A(flit222[5]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][5]));
	BUFX1 U1931(.A(flit222[6]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][6]));
	BUFX1 U1932(.A(flit222[7]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][7]));
	BUFX1 U1933(.A(flit222[8]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][8]));
	BUFX1 U1934(.A(flit222[9]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][9]));
	BUFX1 U1935(.A(flit222[10]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][10]));
	BUFX1 U1936(.A(flit222[11]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][11]));
	BUFX1 U1937(.A(flit222[12]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][12]));
	BUFX1 U1938(.A(flit222[13]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][13]));
	BUFX1 U1939(.A(flit222[14]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][14]));
	BUFX1 U1940(.A(flit222[15]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][15]));
	BUFX1 U1941(.A(flit222[16]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][16]));
	BUFX1 U1942(.A(flit222[17]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][17]));
	BUFX1 U1943(.A(flit222[18]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][18]));
	BUFX1 U1944(.A(flit222[19]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][19]));
	BUFX1 U1945(.A(flit222[20]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][20]));
	BUFX1 U1946(.A(flit222[21]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][21]));
	BUFX1 U1947(.A(flit222[22]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][22]));
	BUFX1 U1948(.A(flit222[23]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][23]));
	BUFX1 U1949(.A(flit222[24]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][24]));
	BUFX1 U1950(.A(flit222[25]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][25]));
	BUFX1 U1951(.A(flit222[26]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][26]));
	BUFX1 U1952(.A(flit222[27]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][27]));
	BUFX1 U1953(.A(flit222[28]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][28]));
	BUFX1 U1954(.A(flit222[29]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][29]));
	BUFX1 U1955(.A(flit222[30]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][30]));
	BUFX1 U1956(.A(flit222[31]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][31]));
	BUFX1 U1957(.A(flit222[32]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][32]));
	BUFX1 U1958(.A(flit222[33]), .Y(from_input_req_in_jump_input_datapath2put_datapath2[110:77][33]));
    NOR2X1 U1959 ( .IN1(flit222[33]), .IN2(flit222[32]), .QN(norres_vc_buffer222_vc_buffer2) );
    OR4X1 U1960 ( .IN1(flit222[29]), .IN2(flit222[28]), .IN3(flit222[27]), .IN4(flit222[26]), .Y(or1res_vc_buffer222) );
    OR4X1 U1961 ( .IN1(flit222[25]), .IN2(flit222[24]), .IN3(flit222[23]), .IN4(flit222[22]), .Y(or2res_vc_buffer222) );
    OR2X1 U1962 ( .A(or1res_vc_buffer222), .B(or2res_vc_buffer222), .Y(orres_vc_buffer222) );
    AND3X1 U1963 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(norres_vc_buffer222_vc_buffer2), .IN3(orres_vc_buffer222), .Q(finres1_vc_buffer222) );
    MUX21X1 U1964 (.IN1(next_locked_vc_buffer222), .IN2(1'b1), .S(finres1_vc_buffer222), .Q(next_locked_vc_buffer222);
    AND3X1 U1965 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(flit222[33]), .IN3(flit222[32]), .Q(andres1_vc_buffer222) );
    MUX21X1 U1966 (.IN1(next_locked_vc_buffer222), .IN2(1'b0), .S(andres1_vc_buffer222), .Q(next_locked_vc_buffer222);

    INVX1 U1967 ( .A(full_vc_buffer222), .Y(full_vc_buffer222_not2) );
    INVX1 U1968 ( .A(locked_by_route_ff_vc_buffer222), .Y(locked_by_route_ff_vc_buffer222_not2) );

    MUX21X1 U1969 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer222_not2), .S(norres_vc_buffer222_vc_buffer2), .Q(thirdand_vc_buffer222);
    AND3X1 U1970 ( .IN1(from_input_req_in_jump_input_datapath2put_datapath2[74]), .IN2(full_vc_buffer222_not2), .IN3(thirdand_vc_buffer222), .Q(write_flit222_vc_buffer22) );
    AND2X1 U1971 ( .IN1(full_vc_buffer222_not2), .IN2(norres_vc_buffer222_vc_buffer2), .Q(from_input_resp_input_datapath2[2]) );
    INVX1 U1972 ( .A(empty_vc_buffer222), .Y(to_output_req_in_jump_input_datapath2put_datapath2[74]) );
    AND2X1 U1973 ( .IN1(to_output_req_in_jump_input_datapath2put_datapath2[74]), .IN2(to_output_resp_input_datapath2[2]), .Q(read_flit222_vc_buffer22) );
	BUFX1 U1974(.A(to_output_req_in_jump_input_datapath2put_datapath2[76:75]), .Y(2'b10));

	DFFX2 U1975 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U1976 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U1977 (.IN1(next_locked_vc_buffer222), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer222);

	BUFX1 U1978(.A(from_input_req_in_jump_input_datapath2put_datapath2[77]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U1979(.A(from_input_req_in_jump_input_datapath2put_datapath2[78]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U1980(.A(from_input_req_in_jump_input_datapath2put_datapath2[79]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U1981(.A(from_input_req_in_jump_input_datapath2put_datapath2[80]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U1982(.A(from_input_req_in_jump_input_datapath2put_datapath2[81]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U1983(.A(from_input_req_in_jump_input_datapath2put_datapath2[82]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U1984(.A(from_input_req_in_jump_input_datapath2put_datapath2[83]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U1985(.A(from_input_req_in_jump_input_datapath2put_datapath2[84]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U1986(.A(from_input_req_in_jump_input_datapath2put_datapath2[85]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U1987(.A(from_input_req_in_jump_input_datapath2put_datapath2[86]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U1988(.A(from_input_req_in_jump_input_datapath2put_datapath2[87]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U1989(.A(from_input_req_in_jump_input_datapath2put_datapath2[88]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U1990(.A(from_input_req_in_jump_input_datapath2put_datapath2[89]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U1991(.A(from_input_req_in_jump_input_datapath2put_datapath2[90]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U1992(.A(from_input_req_in_jump_input_datapath2put_datapath2[91]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U1993(.A(from_input_req_in_jump_input_datapath2put_datapath2[92]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U1994(.A(from_input_req_in_jump_input_datapath2put_datapath2[93]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U1995(.A(from_input_req_in_jump_input_datapath2put_datapath2[94]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U1996(.A(from_input_req_in_jump_input_datapath2put_datapath2[95]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U1997(.A(from_input_req_in_jump_input_datapath2put_datapath2[96]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U1998(.A(from_input_req_in_jump_input_datapath2put_datapath2[97]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U1999(.A(from_input_req_in_jump_input_datapath2put_datapath2[98]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U2000(.A(from_input_req_in_jump_input_datapath2put_datapath2[99]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U2001(.A(from_input_req_in_jump_input_datapath2put_datapath2[100]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U2002(.A(from_input_req_in_jump_input_datapath2put_datapath2[101]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U2003(.A(from_input_req_in_jump_input_datapath2put_datapath2[102]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U2004(.A(from_input_req_in_jump_input_datapath2put_datapath2[103]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U2005(.A(from_input_req_in_jump_input_datapath2put_datapath2[104]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U2006(.A(from_input_req_in_jump_input_datapath2put_datapath2[105]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U2007(.A(from_input_req_in_jump_input_datapath2put_datapath2[106]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U2008(.A(from_input_req_in_jump_input_datapath2put_datapath2[107]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U2009(.A(from_input_req_in_jump_input_datapath2put_datapath2[108]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U2010(.A(from_input_req_in_jump_input_datapath2put_datapath2[109]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U2011(.A(from_input_req_in_jump_input_datapath2put_datapath2[110]), .Y(ext_req_v_i[110:74][36]));
    XNOR2X1 U2012 ( .IN1(ext_req_v_i[110:74][1]), .IN2(i_input_datapath2[0]), .QN(xnor1resu_input_datapath2) );
    XNOR2X1 U2013 ( .IN1(ext_req_v_i[110:74][2]), .IN2(i_input_datapath2[1]), .QN(xnor2resu_input_datapath2) );
    AND2X1 U2014 ( .IN1(xnor1resu_input_datapath2), .IN2(xnor2resu_input_datapath2), .Q(and1resu_input_datapath2) );
    AND3X1 U2015 ( .IN1(and1resu_input_datapath2), .IN2(ext_req_v_i[110:74][0]), .IN2(ext_req_v_i[110:74][0]), .Q(cond1line_input_datapath2) );
    MUX21X1 U2016 (.IN1(vc_ch_act_in_input_datapath2[0]), .IN2(i_input_datapath2[0]), .S(cond1line_input_datapath2), .Q(vc_ch_act_in_input_datapath2[0]));
    MUX21X1 U2017 (.IN1(vc_ch_act_in_input_datapath2[1]), .IN2(i_input_datapath2[1]), .S(cond1line_input_datapath2), .Q(vc_ch_act_in_input_datapath2[1]));
    MUX21X1 U2018 (.IN1(req_in_jump_input_datapath2), .IN2(1), .S(cond1line_input_datapath2), .Q(req_in_jump_input_datapath2));
	BUFX1 U2019(.A(from_input_req_in_jump_input_datapath2put_datapath2[40]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U2020(.A(from_input_req_in_jump_input_datapath2put_datapath2[41]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U2021(.A(from_input_req_in_jump_input_datapath2put_datapath2[42]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U2022(.A(from_input_req_in_jump_input_datapath2put_datapath2[43]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U2023(.A(from_input_req_in_jump_input_datapath2put_datapath2[44]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U2024(.A(from_input_req_in_jump_input_datapath2put_datapath2[45]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U2025(.A(from_input_req_in_jump_input_datapath2put_datapath2[46]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U2026(.A(from_input_req_in_jump_input_datapath2put_datapath2[47]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U2027(.A(from_input_req_in_jump_input_datapath2put_datapath2[48]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U2028(.A(from_input_req_in_jump_input_datapath2put_datapath2[49]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U2029(.A(from_input_req_in_jump_input_datapath2put_datapath2[50]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U2030(.A(from_input_req_in_jump_input_datapath2put_datapath2[51]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U2031(.A(from_input_req_in_jump_input_datapath2put_datapath2[52]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U2032(.A(from_input_req_in_jump_input_datapath2put_datapath2[53]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U2033(.A(from_input_req_in_jump_input_datapath2put_datapath2[54]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U2034(.A(from_input_req_in_jump_input_datapath2put_datapath2[55]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U2035(.A(from_input_req_in_jump_input_datapath2put_datapath2[56]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U2036(.A(from_input_req_in_jump_input_datapath2put_datapath2[57]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U2037(.A(from_input_req_in_jump_input_datapath2put_datapath2[58]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U2038(.A(from_input_req_in_jump_input_datapath2put_datapath2[59]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U2039(.A(from_input_req_in_jump_input_datapath2put_datapath2[60]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U2040(.A(from_input_req_in_jump_input_datapath2put_datapath2[61]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U2041(.A(from_input_req_in_jump_input_datapath2put_datapath2[62]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U2042(.A(from_input_req_in_jump_input_datapath2put_datapath2[63]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U2043(.A(from_input_req_in_jump_input_datapath2put_datapath2[64]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U2044(.A(from_input_req_in_jump_input_datapath2put_datapath2[65]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U2045(.A(from_input_req_in_jump_input_datapath2put_datapath2[66]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U2046(.A(from_input_req_in_jump_input_datapath2put_datapath2[67]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U2047(.A(from_input_req_in_jump_input_datapath2put_datapath2[68]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U2048(.A(from_input_req_in_jump_input_datapath2put_datapath2[69]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U2049(.A(from_input_req_in_jump_input_datapath2put_datapath2[70]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U2050(.A(from_input_req_in_jump_input_datapath2put_datapath2[71]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U2051(.A(from_input_req_in_jump_input_datapath2put_datapath2[72]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U2052(.A(from_input_req_in_jump_input_datapath2put_datapath2[73]), .Y(ext_req_v_i[110:74][36]));

	BUFX1 U2053(.A(from_input_req_in_jump_input_datapath2put_datapath2[3]), .Y(ext_req_v_i[110:74][3]));
	BUFX1 U2054(.A(from_input_req_in_jump_input_datapath2put_datapath2[4]), .Y(ext_req_v_i[110:74][4]));
	BUFX1 U2055(.A(from_input_req_in_jump_input_datapath2put_datapath2[5]), .Y(ext_req_v_i[110:74][5]));
	BUFX1 U2056(.A(from_input_req_in_jump_input_datapath2put_datapath2[6]), .Y(ext_req_v_i[110:74][6]));
	BUFX1 U2057(.A(from_input_req_in_jump_input_datapath2put_datapath2[7]), .Y(ext_req_v_i[110:74][7]));
	BUFX1 U2058(.A(from_input_req_in_jump_input_datapath2put_datapath2[8]), .Y(ext_req_v_i[110:74][8]));
	BUFX1 U2059(.A(from_input_req_in_jump_input_datapath2put_datapath2[9]), .Y(ext_req_v_i[110:74][9]));
	BUFX1 U2060(.A(from_input_req_in_jump_input_datapath2put_datapath2[10]), .Y(ext_req_v_i[110:74][10]));
	BUFX1 U2061(.A(from_input_req_in_jump_input_datapath2put_datapath2[11]), .Y(ext_req_v_i[110:74][11]));
	BUFX1 U2062(.A(from_input_req_in_jump_input_datapath2put_datapath2[12]), .Y(ext_req_v_i[110:74][12]));
	BUFX1 U2063(.A(from_input_req_in_jump_input_datapath2put_datapath2[13]), .Y(ext_req_v_i[110:74][13]));
	BUFX1 U2064(.A(from_input_req_in_jump_input_datapath2put_datapath2[14]), .Y(ext_req_v_i[110:74][14]));
	BUFX1 U2065(.A(from_input_req_in_jump_input_datapath2put_datapath2[15]), .Y(ext_req_v_i[110:74][15]));
	BUFX1 U2066(.A(from_input_req_in_jump_input_datapath2put_datapath2[16]), .Y(ext_req_v_i[110:74][16]));
	BUFX1 U2067(.A(from_input_req_in_jump_input_datapath2put_datapath2[17]), .Y(ext_req_v_i[110:74][17]));
	BUFX1 U2068(.A(from_input_req_in_jump_input_datapath2put_datapath2[18]), .Y(ext_req_v_i[110:74][18]));
	BUFX1 U2069(.A(from_input_req_in_jump_input_datapath2put_datapath2[19]), .Y(ext_req_v_i[110:74][19]));
	BUFX1 U2070(.A(from_input_req_in_jump_input_datapath2put_datapath2[20]), .Y(ext_req_v_i[110:74][20]));
	BUFX1 U2071(.A(from_input_req_in_jump_input_datapath2put_datapath2[21]), .Y(ext_req_v_i[110:74][21]));
	BUFX1 U2072(.A(from_input_req_in_jump_input_datapath2put_datapath2[22]), .Y(ext_req_v_i[110:74][22]));
	BUFX1 U2073(.A(from_input_req_in_jump_input_datapath2put_datapath2[23]), .Y(ext_req_v_i[110:74][23]));
	BUFX1 U2074(.A(from_input_req_in_jump_input_datapath2put_datapath2[24]), .Y(ext_req_v_i[110:74][24]));
	BUFX1 U2075(.A(from_input_req_in_jump_input_datapath2put_datapath2[25]), .Y(ext_req_v_i[110:74][25]));
	BUFX1 U2076(.A(from_input_req_in_jump_input_datapath2put_datapath2[26]), .Y(ext_req_v_i[110:74][26]));
	BUFX1 U2077(.A(from_input_req_in_jump_input_datapath2put_datapath2[27]), .Y(ext_req_v_i[110:74][27]));
	BUFX1 U2078(.A(from_input_req_in_jump_input_datapath2put_datapath2[28]), .Y(ext_req_v_i[110:74][28]));
	BUFX1 U2079(.A(from_input_req_in_jump_input_datapath2put_datapath2[29]), .Y(ext_req_v_i[110:74][29]));
	BUFX1 U2080(.A(from_input_req_in_jump_input_datapath2put_datapath2[30]), .Y(ext_req_v_i[110:74][30]));
	BUFX1 U2081(.A(from_input_req_in_jump_input_datapath2put_datapath2[31]), .Y(ext_req_v_i[110:74][31]));
	BUFX1 U2082(.A(from_input_req_in_jump_input_datapath2put_datapath2[32]), .Y(ext_req_v_i[110:74][32]));
	BUFX1 U2083(.A(from_input_req_in_jump_input_datapath2put_datapath2[33]), .Y(ext_req_v_i[110:74][33]));
	BUFX1 U2084(.A(from_input_req_in_jump_input_datapath2put_datapath2[34]), .Y(ext_req_v_i[110:74][34]));
	BUFX1 U2085(.A(from_input_req_in_jump_input_datapath2put_datapath2[35]), .Y(ext_req_v_i[110:74][35]));
	BUFX1 U2086(.A(from_input_req_in_jump_input_datapath2put_datapath2[36]), .Y(ext_req_v_i[110:74][36]));

    MUX21X1 U2087 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2 * 37]), .IN2(ext_req_v_i[110:74][0]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2 * 37]));
    MUX21X1 U2088 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+2]), .IN2(vc_ch_act_in_input_datapath2[1]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+2]));
    MUX21X1 U2089 (.IN1(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+1]), .IN2(vc_ch_act_in_input_datapath2[0]), .S(req_in_jump_input_datapath2), .Q(from_input_req_in_jump_input_datapath2put_datapath2[vc_ch_act_in_input_datapath2*37+1]));
    MUX21X1 U2090 (.IN1(ext_resp_v_o[3:2][0]), .IN2(from_input_resp_input_datapath2[vc_ch_act_in_input_datapath2]), .S(req_in_jump_input_datapath2), .Q(ext_resp_v_o[3:2][0]));

    INVX1 U2091 ( .A(req_in_jump_input_datapath2), .Y(req_in_jump_input_datapath2_not) );
    MUX21X1 U2092 (.IN1(ext_resp_v_o[3:2][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath2_not), .Q(ext_resp_v_o[3:2][0]));
    BUFX1 U2093(.A(from_input_req_in_jump_input_datapath2put_datapath2[34]), .Y(ext_req_v_i[110:74][34]));

    XOR2X1 U2094 ( .IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b1), .Q(xor1resu_input_datapath2) );
    MUX21X1 U2095 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(xor1resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U2096 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b0), .S(xor1resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[1]));
    AND2X1 U2097 ( .IN1(xor1resu_input_datapath2), .IN2(to_output_req_in_jump_input_datapath2put_datapath2[j_input_datapath2*37]), .Q(and2resu_input_datapath2) );
    MUX21X1 U2098 (.IN1(vc_ch_act_out_input_datapath2[0]), .IN2(j_input_datapath2[0]), .S(and2resu_input_datapath2), .Q(vc_ch_act_out_input_datapath2[0]));
    MUX21X1 U2099 (.IN1(vc_ch_act_out_input_datapath2[1]), .IN2(j_input_datapath2[1]), .S(and2resu_input_datapath2), .Q(vc_ch_act_out_input_datapath2[1]));
    MUX21X1 U2100 (.IN1(req_out_jump_input_datapath2), .IN2(1'b1), .S(and2resu_input_datapath2), .Q(req_out_jump_input_datapath2));
    MUX21X1 U2101 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(and2resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U2102 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b1), .S(and2resu_input_datapath2), .Q(_sv2v_jump_input_datapath2[1]));
    HADDX1 U2103 ( .A0(j_input_datapath2[0]), .B0(1'b1), .C1(j_input_datapath2[1]), .SO(j_input_datapath2[0]) );
    HADDX1 U2104 ( .A0(j_input_datapath2[0]), .B0(1'b1), .C1(j_input_datapath2[1]), .SO(j_input_datapath2[0]) );
    AND2X1 U2105 ( .IN1(xor1resu_input_datapath2), .IN2(to_output_req_in_jump_input_datapath2put_datapath2[j_input_datapath2*37]), .Q(and3resu) );
    NAND2X1 U2106(.A(_sv2v_jump_input_datapath2[0]),.B(_sv2v_jump_input_datapath2[1]),.Y(nand1resu_input_datapath22));
    MUX21X1 U2107 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(1'b0), .S(nand1resu_input_datapath22), .Q(_sv2v_jump_input_datapath2[0]));
    MUX21X1 U2108 (.IN1(_sv2v_jump_input_datapath2[1]), .IN2(1'b0), .S(nand1resu_input_datapath22), .Q(_sv2v_jump_input_datapath2[1]));
    XNOR2X1 U2109 (.IN1(_sv2v_jump_input_datapath2[0]), .IN2(_sv2v_jump_input_datapath2[1]), .Q(xnor23resu_input_datapath2) );
    AND2X1 U2110 ( .IN1(xnor23resu_input_datapath2), .IN2(req_out_jump_input_datapath2), .Q(and4resu_input_datapath2) );

    MUX21X1 U2111(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[110:74][3]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U2112(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[110:74][4]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U2113(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[110:74][5]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U2114(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[110:74][6]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U2115(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[110:74][7]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U2116(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[110:74][8]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U2117(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[110:74][9]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U2118(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[110:74][10]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U2119(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[110:74][11]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U2120(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[110:74][12]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U2121(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[110:74][13]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U2122(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[110:74][14]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U2123(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[110:74][15]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U2124(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[110:74][16]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U2125(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[110:74][17]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U2126(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[110:74][18]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U2127(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[110:74][19]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U2128(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[110:74][20]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U2129(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[110:74][21]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U2130(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[110:74][22]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U2131(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[110:74][23]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U2132(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[110:74][24]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U2133(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[110:74][25]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U2134(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[110:74][26]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U2135(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[110:74][27]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U2136(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[110:74][28]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U2137(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[110:74][29]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U2138(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[110:74][30]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U2139(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[110:74][31]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U2140(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[110:74][32]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U2141(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[110:74][33]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U2142(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[110:74][34]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U2143(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[110:74][35]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U2144(.IN1(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[110:74][36]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U2145(.IN1(int_req_v[110:74][0]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2 * 37)]), .S(and4resu_input_datapath2), .Q(int_req_v[110:74][0]));
	MUX21X1 U2146(.IN1(int_req_v[110:74][1]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+1]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+1]));
	MUX21X1 U2147(.IN1(int_req_v[110:74][2]),.IN2(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+2]), .S(and4resu_input_datapath2), .Q(to_output_req_in_jump_input_datapath2put_datapath2[(vc_ch_act_out_input_datapath2*37)+2]));
	MUX21X1 U2148(.IN1(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2]),.IN2(int_resp_v[3:2]), .S(and4resu_input_datapath2), .Q(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2]));
	MUX21X1 U2149(.IN1(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2+1]),.IN2(int_resp_v[3:2]), .S(and4resu_input_datapath2), .Q(to_output_resp_input_datapath2[vc_ch_act_out_input_datapath2+1]));


	BUFX1 U2150 ( .A(read_ptr_ff_fifomodule3[0]), .Y(next_read_ptr_fifomodule3[0]) );
	BUFX1 U2151 ( .A(read_ptr_ff_fifomodule3[1]), .Y(next_read_ptr_fifomodule3[1]) );
	BUFX1 U2152 ( .A(write_ptr_ff_fifomodule3[0]), .Y(next_write_ptr_fifomodule3[0]) );
	BUFX1 U2153 ( .A(write_ptr_ff_fifomodule3[1]), .Y(next_write_ptr_fifomodule3[1]) );

	XNOR2X1 U2154 ( .IN1(write_ptr_ff_fifomodule3[0]), .IN2(read_ptr_ff_fifomodule3[0]), .Q(u1temp_fifomodule3) );
	XNOR2X1 U2155 ( .IN1(write_ptr_ff_fifomodule3[1]), .IN2(read_ptr_ff_fifomodule3[1]), .Q(u2temp_fifomodule3) );
	AND2X1 U2156 ( .A(u1temp_fifomodule3), .B(u2temp_fifomodule3), .Y(empty_vc_buffer3) );
	XOR2X1 U2157 ( .A(write_ptr_ff_fifomodule3[1]), .B(read_ptr_ff_fifomodule3[1]), .Y(u4temp_fifomodule3) );
	AND2X1 U2158 ( .A(u1temp_fifomodule3), .B(u4temp_fifomodule3), .Y(full_vc_buffer3) );
	MUX21X1 U2159 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][0]));
	MUX21X1 U2160 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][1]));
	MUX21X1 U2161 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][2]));
	MUX21X1 U2162 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][3]));
	MUX21X1 U2163 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][4]));
	MUX21X1 U2164 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][5]));
	MUX21X1 U2165 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][6]));
	MUX21X1 U2166 (.IN1(fifo_ff_fifomodule3[read_ptr_ff_fifomodule3[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[36:3][7]));

	INVX1 U2167 ( .A(full_vc_buffer3), .Y(full_vc_buffer3_not_fifomodule) );
	AND2X1 U2168 ( .A(write_flit3_vc_buffer3), .B(full_vc_buffer3_not_fifomodule), .Y(u7temp_fifomodule3) );
	MUX21X1 U2169 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule3), .Q(u9temp_fifomodule3));
	HADDX1 U2170 ( .A0(write_ptr_ff_fifomodule3[0]), .B0(u9temp_fifomodule3), .C1(u10carry_fifomodule3), .SO(next_write_ptr_fifomodule3[0]) );
	HADDX1 U2171 ( .A0(u10carry_fifomodule3), .B0(write_ptr_ff_fifomodule3[1]), .C1(u11carry_fifomodule3), .SO(next_write_ptr_fifomodule3[1]) );

	INVX1 U2172 ( .A(empty_vc_buffer3), .Y(empty_vc_buffer3_not_fifomodule) );
	AND2X1 U2173 ( .A(read_flit3_vc_buffer3), .B(empty_vc_buffer3_not_fifomodule), .Y(u13temp_fifomodule3) );
	MUX21X1 U2174 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule3), .Q(u14temp_fifomodule3));
	HADDX1 U2175 ( .A0(read_ptr_ff_fifomodule3[0]), .B0(u14temp_fifomodule3), .C1(u15carry_fifomodule3), .SO(next_read_ptr_fifomodule3[0]) );
	HADDX1 U2176 ( .A0(u15carry_fifomodule3), .B0(read_ptr_ff_fifomodule3[1]), .C1(u16carry_fifomodule3), .SO(next_read_ptr_fifomodule3[1]) );

	AND2X1 U2177 ( .A(write_flit3_vc_buffer3), .B(full_vc_buffer3), .Y(u17res_fifomodule3) );
	AND2X1 U2178 ( .A(read_flit3_vc_buffer3), .B(empty_vc_buffer3), .Y(u18res_fifomodule3) );
    OR2X1 U2179 ( .A(u17res_fifomodule3), .B(u18res_fifomodule3), .Y(error_vc_buffer3) );
	XOR2X1 U2180 ( .A(write_ptr_ff_fifomodule3[0]), .B(read_ptr_ff_fifomodule3[0]), .Y(fifo_ocup_fifomodule3[0]) );
	INVX1 U2181 ( .A(write_ptr_ff_fifomodule3[0]), .Y(write_ptr_ff_fifomodule3_0_not3) );
	AND2X1 U2182 ( .A(write_ptr_ff_fifomodule3_0_not3), .B(read_ptr_ff_fifomodule3[0]), .Y(b0wire_fifomodule3) );
	XOR2X1 U2183 ( .A(write_ptr_ff_fifomodule3[1]), .B(read_ptr_ff_fifomodule3[1]), .Y(u23temp_fifomodule3) );
	INVX1 U2184 ( .A(write_ptr_ff_fifomodule3[1]), .Y(write_ptr_ff_fifomodule3_1_not3) );
	AND2X1 U2185 ( .A(read_ptr_ff_fifomodule3[1]), .B(write_ptr_ff_fifomodule3_1_not3), .Y(boutb_fifomodule3) );
	XOR2X1 U2186 ( .A(u23temp_fifomodule3), .B(b0wire_fifomodule3), .Y(fifo_ocup_fifomodule3[1]) );
	INVX1 U2187 ( .A(u23temp_fifomodule3), .Y(u23temp_fifomodule3_not_fifomodule3) );
	AND2X1 U2188 ( .A(b0wire_fifomodule3), .B(u23temp_fifomodule3_not_fifomodule3), .Y(bouta_fifomodule3) );
	OR2X1 U2189 ( .A(bouta_fifomodule3), .B(boutb_fifomodule3), .Y(boutmain_fifomodule3) );
	DFFX2 U2190 ( .CLK(clk), .D(fifo_ocup_fifomodule3[0]), .Q(ocup_o[0]) );
	DFFX2 U2191 ( .CLK(clk), .D(fifo_ocup_fifomodule3[1]), .Q(ocup_o[1]) );
	DFFX2 U2192 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule3) );
	DFFX2 U2193 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule3) );
	DFFX2 U2194 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(write_ptr_ff_fifomodule3[0]) );
	DFFX2 U2195 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(read_ptr_ff_fifomodule3[0]) );
	DFFX2 U2196 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(fifo_ff_fifomodule3[0]) );
	DFFX2 U2197 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(write_ptr_ff_fifomodule3[1]) );
	DFFX2 U2198 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(read_ptr_ff_fifomodule3[1]) );
	DFFX2 U2199 ( .CLK(arst_value_fifomodule3), .D(1'b0), .Q(fifo_ff_fifomodule3[1]) );

	DFFX2 U2200 ( .CLK(clk), .D(next_write_ptr_fifomodule3[0]), .Q(write_ptr_ff_fifomodule3[0]) );
	DFFX2 U2201 ( .CLK(clk), .D(next_write_ptr_fifomodule3[1]), .Q(write_ptr_ff_fifomodule3[1]) );
	DFFX2 U2202 ( .CLK(clk), .D(next_read_ptr_fifomodule3[0]), .Q(read_ptr_ff_fifomodule3[0]) );
	DFFX2 U2203 ( .CLK(clk), .D(next_read_ptr_fifomodule3[1]), .Q(read_ptr_ff_fifomodule3[1]) );
	  

	DFFX2 U2204 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][0]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8]) );
	DFFX2 U2205 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][1]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+1]) );
	DFFX2 U2206 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][2]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+2]) );
	DFFX2 U2207 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][3]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+3]) );
	DFFX2 U2208 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][4]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+4]) );
	DFFX2 U2209 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][5]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+5]) );
	DFFX2 U2210 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][6]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+6]) );
	DFFX2 U2211 ( .CLK(u7temp_fifomodule3), .D(from_input_req_in_jump_input_datapath3put_datapath3[36:3][7]), .Q(fifo_ff_fifomodule3[write_ptr_ff_fifomodule3[0]*8+7]) );

    BUFX1 U2212 ( .A(locked_by_route_ff_vc_buffer3), .Y(next_locked_vc_buffer3) );
    BUFX1 U2213(.A(flit3[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][0]));
	BUFX1 U2214(.A(flit3[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][1]));
	BUFX1 U2215(.A(flit3[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][2]));
	BUFX1 U2216(.A(flit3[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][3]));
	BUFX1 U2217(.A(flit3[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][4]));
	BUFX1 U2218(.A(flit3[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][5]));
	BUFX1 U2219(.A(flit3[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][6]));
	BUFX1 U2220(.A(flit3[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][7]));
	BUFX1 U2221(.A(flit3[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][8]));
	BUFX1 U2222(.A(flit3[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][9]));
	BUFX1 U2223(.A(flit3[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][10]));
	BUFX1 U2224(.A(flit3[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][11]));
	BUFX1 U2225(.A(flit3[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][12]));
	BUFX1 U2226(.A(flit3[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][13]));
	BUFX1 U2227(.A(flit3[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][14]));
	BUFX1 U2228(.A(flit3[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][15]));
	BUFX1 U2229(.A(flit3[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][16]));
	BUFX1 U2230(.A(flit3[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][17]));
	BUFX1 U2231(.A(flit3[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][18]));
	BUFX1 U2232(.A(flit3[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][19]));
	BUFX1 U2233(.A(flit3[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][20]));
	BUFX1 U2234(.A(flit3[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][21]));
	BUFX1 U2235(.A(flit3[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][22]));
	BUFX1 U2236(.A(flit3[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][23]));
	BUFX1 U2237(.A(flit3[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][24]));
	BUFX1 U2238(.A(flit3[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][25]));
	BUFX1 U2239(.A(flit3[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][26]));
	BUFX1 U2240(.A(flit3[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][27]));
	BUFX1 U2241(.A(flit3[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][28]));
	BUFX1 U2242(.A(flit3[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][29]));
	BUFX1 U2243(.A(flit3[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][30]));
	BUFX1 U2244(.A(flit3[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][31]));
	BUFX1 U2245(.A(flit3[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][32]));
	BUFX1 U2246(.A(flit3[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[36:3][33]));
    NOR2X1 U2247 ( .IN1(flit3[33]), .IN2(flit3[32]), .QN(norres_vc_buffer3_vc_buffer3) );
    OR4X1 U2248 ( .IN1(flit3[29]), .IN2(flit3[28]), .IN3(flit3[27]), .IN4(flit3[26]), .Y(or1res_vc_buffer3) );
    OR4X1 U2249 ( .IN1(flit3[25]), .IN2(flit3[24]), .IN3(flit3[23]), .IN4(flit3[22]), .Y(or2res_vc_buffer3) );
    OR2X1 U2250 ( .A(or1res_vc_buffer3), .B(or2res_vc_buffer3), .Y(orres_vc_buffer3) );
    AND3X1 U2251 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(norres_vc_buffer3_vc_buffer3), .IN3(orres_vc_buffer3), .Q(finres1_vc_buffer3) );
    MUX21X1 U2252 (.IN1(next_locked_vc_buffer3), .IN2(1'b1), .S(finres1_vc_buffer3), .Q(next_locked_vc_buffer3);
    AND3X1 U2253 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(flit3[33]), .IN3(flit3[32]), .Q(andres1_vc_buffer3) );
    MUX21X1 U2254 (.IN1(next_locked_vc_buffer3), .IN2(1'b0), .S(andres1_vc_buffer3), .Q(next_locked_vc_buffer3);

    INVX1 U2255 ( .A(full_vc_buffer3), .Y(full_vc_buffer3_not) );
    INVX1 U2256 ( .A(locked_by_route_ff_vc_buffer3), .Y(locked_by_route_ff_vc_buffer3_not) );

    MUX21X1 U2257 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer3_not), .S(norres_vc_buffer3_vc_buffer3), .Q(thirdand_vc_buffer3);
    AND3X1 U2258 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[0]), .IN2(full_vc_buffer3_not), .IN3(thirdand_vc_buffer3), .Q(write_flit3_vc_buffer3) );
    AND2X1 U2259 ( .IN1(full_vc_buffer3_not), .IN2(norres_vc_buffer3_vc_buffer3), .Q(from_input_resp_input_datapath3[0]) );
    INVX1 U2260 ( .A(empty_vc_buffer3), .Y(to_output_req_in_jump_input_datapath3put_datapath3[0]) );
    AND2X1 U2261 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[0]), .IN2(to_output_resp_input_datapath3[0]), .Q(read_flit3_vc_buffer3) );
	BUFX1 U2262(.A(to_output_req_in_jump_input_datapath3put_datapath3[2:1]), .Y(2'b00));

	DFFX2 U2263 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U2264 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U2265 (.IN1(next_locked_vc_buffer3), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer3);

	BUFX1 U2266 ( .A(read_ptr_ff_fifomodule31[0]), .Y(next_read_ptr_fifomodule31[0]) );
	BUFX1 U2267 ( .A(read_ptr_ff_fifomodule31[1]), .Y(next_read_ptr_fifomodule31[1]) );
	BUFX1 U2268 ( .A(write_ptr_ff_fifomodule31[0]), .Y(next_write_ptr_fifomodule31[0]) );
	BUFX1 U2269 ( .A(write_ptr_ff_fifomodule31[1]), .Y(next_write_ptr_fifomodule31[1]) );

	XNOR2X1 U2270 ( .IN1(write_ptr_ff_fifomodule31[0]), .IN2(read_ptr_ff_fifomodule31[0]), .Q(u1temp_fifomodule31) );
	XNOR2X1 U2271 ( .IN1(write_ptr_ff_fifomodule31[1]), .IN2(read_ptr_ff_fifomodule31[1]), .Q(u2temp_fifomodule31) );
	AND2X1 U2272 ( .A(u1temp_fifomodule31), .B(u2temp_fifomodule31), .Y(empty_vc_buffer31) );
	XOR2X1 U2273 ( .A(write_ptr_ff_fifomodule31[1]), .B(read_ptr_ff_fifomodule31[1]), .Y(u4temp_fifomodule31) );
	AND2X1 U2274 ( .A(u1temp_fifomodule31), .B(u4temp_fifomodule31), .Y(full_vc_buffer31) );
	MUX21X1 U2275 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][0]));
	MUX21X1 U2276 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][1]));
	MUX21X1 U2277 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][2]));
	MUX21X1 U2278 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][3]));
	MUX21X1 U2279 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][4]));
	MUX21X1 U2280 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][5]));
	MUX21X1 U2281 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][6]));
	MUX21X1 U2282 (.IN1(fifo_ff_fifomodule31[read_ptr_ff_fifomodule31[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer31), .Q(to_output_req_in_jump_input_datapath3put_datapath3[73:40][7]));

	INVX1 U2283 ( .A(full_vc_buffer31), .Y(full_vc_buffer31_not1_fifomodule1) );
	AND2X1 U2284 ( .A(write_flit31_vc_buffer13), .B(full_vc_buffer31_not1_fifomodule1), .Y(u7temp_fifomodule31) );
	MUX21X1 U2285 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule31), .Q(u9temp_fifomodule31));
	HADDX1 U2286 ( .A0(write_ptr_ff_fifomodule31[0]), .B0(u9temp_fifomodule31), .C1(u10carry_fifomodule31), .SO(next_write_ptr_fifomodule31[0]) );
	HADDX1 U2287 ( .A0(u10carry_fifomodule31), .B0(write_ptr_ff_fifomodule31[1]), .C1(u11carry_fifomodule31), .SO(next_write_ptr_fifomodule31[1]) );

	INVX1 U2288 ( .A(empty_vc_buffer31), .Y(empty_vc_buffer31_not_fifomodule1) );
	AND2X1 U2289 ( .A(read_flit31_vc_buffer13), .B(empty_vc_buffer31_not_fifomodule1), .Y(u13temp_fifomodule31) );
	MUX21X1 U2290 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule31), .Q(u14temp_fifomodule31));
	HADDX1 U2291 ( .A0(read_ptr_ff_fifomodule31[0]), .B0(u14temp_fifomodule31), .C1(u15carry_fifomodule31), .SO(next_read_ptr_fifomodule31[0]) );
	HADDX1 U2292 ( .A0(u15carry_fifomodule31), .B0(read_ptr_ff_fifomodule31[1]), .C1(u16carry_fifomodule31), .SO(next_read_ptr_fifomodule31[1]) );

	AND2X1 U2293 ( .A(write_flit31_vc_buffer13), .B(full_vc_buffer31), .Y(u17res_fifomodule31) );
	AND2X1 U2294 ( .A(read_flit31_vc_buffer13), .B(empty_vc_buffer31), .Y(u18res_fifomodule31) );
    OR2X1 U2295 ( .A(u17res_fifomodule31), .B(u18res_fifomodule31), .Y(error_vc_buffer31) );
	XOR2X1 U2296 ( .A(write_ptr_ff_fifomodule31[0]), .B(read_ptr_ff_fifomodule31[0]), .Y(fifo_ocup_fifomodule31[0]) );
	INVX1 U2297 ( .A(write_ptr_ff_fifomodule31[0]), .Y(write_ptr_ff_fifomodule31_0_not13) );
	AND2X1 U2298 ( .A(write_ptr_ff_fifomodule31_0_not13), .B(read_ptr_ff_fifomodule31[0]), .Y(b0wire_fifomodule31) );
	XOR2X1 U2299 ( .A(write_ptr_ff_fifomodule31[1]), .B(read_ptr_ff_fifomodule31[1]), .Y(u23temp_fifomodule31) );
	INVX1 U2300 ( .A(write_ptr_ff_fifomodule31[1]), .Y(write_ptr_ff_fifomodule31_1_not13) );
	AND2X1 U2301 ( .A(read_ptr_ff_fifomodule31[1]), .B(write_ptr_ff_fifomodule31_1_not13), .Y(boutb_fifomodule31) );
	XOR2X1 U2302 ( .A(u23temp_fifomodule31), .B(b0wire_fifomodule31), .Y(fifo_ocup_fifomodule31[1]) );
	INVX1 U2303 ( .A(u23temp_fifomodule31), .Y(u23temp_fifomodule31_not_fifomodule1) );
	AND2X1 U2304 ( .A(b0wire_fifomodule31), .B(u23temp_fifomodule31_not_fifomodule1), .Y(bouta_fifomodule31) );
	OR2X1 U2305 ( .A(bouta_fifomodule31), .B(boutb_fifomodule31), .Y(boutmain_fifomodule31) );
	DFFX2 U2306 ( .CLK(clk), .D(fifo_ocup_fifomodule31[0]), .Q(ocup_o[0]) );
	DFFX2 U2307 ( .CLK(clk), .D(fifo_ocup_fifomodule31[1]), .Q(ocup_o[1]) );
	DFFX2 U2308 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule31) );
	DFFX2 U2309 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule31) );
	DFFX2 U2310 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(write_ptr_ff_fifomodule31[0]) );
	DFFX2 U2311 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(read_ptr_ff_fifomodule31[0]) );
	DFFX2 U2312 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(fifo_ff_fifomodule31[0]) );
	DFFX2 U2313 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(write_ptr_ff_fifomodule31[1]) );
	DFFX2 U2314 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(read_ptr_ff_fifomodule31[1]) );
	DFFX2 U2315 ( .CLK(arst_value_fifomodule31), .D(1'b0), .Q(fifo_ff_fifomodule31[1]) );

	DFFX2 U2316 ( .CLK(clk), .D(next_write_ptr_fifomodule31[0]), .Q(write_ptr_ff_fifomodule31[0]) );
	DFFX2 U2317 ( .CLK(clk), .D(next_write_ptr_fifomodule31[1]), .Q(write_ptr_ff_fifomodule31[1]) );
	DFFX2 U2318 ( .CLK(clk), .D(next_read_ptr_fifomodule31[0]), .Q(read_ptr_ff_fifomodule31[0]) );
	DFFX2 U2319 ( .CLK(clk), .D(next_read_ptr_fifomodule31[1]), .Q(read_ptr_ff_fifomodule31[1]) );
	  

	DFFX2 U2320 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][0]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8]) );
	DFFX2 U2321 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][1]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+1]) );
	DFFX2 U2322 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][2]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+2]) );
	DFFX2 U2323 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][3]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+3]) );
	DFFX2 U2324 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][4]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+4]) );
	DFFX2 U2325 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][5]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+5]) );
	DFFX2 U2326 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][6]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+6]) );
	DFFX2 U2327 ( .CLK(u7temp_fifomodule31), .D(from_input_req_in_jump_input_datapath3put_datapath3[73:40][7]), .Q(fifo_ff_fifomodule31[write_ptr_ff_fifomodule31[0]*8+7]) );

    BUFX1 U2328 ( .A(locked_by_route_ff_vc_buffer31), .Y(next_locked_vc_buffer31) );
    BUFX1 U2329(.A(flit31[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][0]));
	BUFX1 U2330(.A(flit31[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][1]));
	BUFX1 U2331(.A(flit31[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][2]));
	BUFX1 U2332(.A(flit31[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][3]));
	BUFX1 U2333(.A(flit31[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][4]));
	BUFX1 U2334(.A(flit31[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][5]));
	BUFX1 U2335(.A(flit31[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][6]));
	BUFX1 U2336(.A(flit31[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][7]));
	BUFX1 U2337(.A(flit31[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][8]));
	BUFX1 U2338(.A(flit31[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][9]));
	BUFX1 U2339(.A(flit31[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][10]));
	BUFX1 U2340(.A(flit31[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][11]));
	BUFX1 U2341(.A(flit31[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][12]));
	BUFX1 U2342(.A(flit31[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][13]));
	BUFX1 U2343(.A(flit31[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][14]));
	BUFX1 U2344(.A(flit31[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][15]));
	BUFX1 U2345(.A(flit31[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][16]));
	BUFX1 U2346(.A(flit31[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][17]));
	BUFX1 U2347(.A(flit31[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][18]));
	BUFX1 U2348(.A(flit31[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][19]));
	BUFX1 U2349(.A(flit31[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][20]));
	BUFX1 U2350(.A(flit31[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][21]));
	BUFX1 U2351(.A(flit31[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][22]));
	BUFX1 U2352(.A(flit31[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][23]));
	BUFX1 U2353(.A(flit31[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][24]));
	BUFX1 U2354(.A(flit31[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][25]));
	BUFX1 U2355(.A(flit31[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][26]));
	BUFX1 U2356(.A(flit31[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][27]));
	BUFX1 U2357(.A(flit31[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][28]));
	BUFX1 U2358(.A(flit31[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][29]));
	BUFX1 U2359(.A(flit31[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][30]));
	BUFX1 U2360(.A(flit31[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][31]));
	BUFX1 U2361(.A(flit31[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][32]));
	BUFX1 U2362(.A(flit31[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[73:40][33]));
    NOR2X1 U2363 ( .IN1(flit31[33]), .IN2(flit31[32]), .QN(norres_vc_buffer31_vc_buffer1) );
    OR4X1 U2364 ( .IN1(flit31[29]), .IN2(flit31[28]), .IN3(flit31[27]), .IN4(flit31[26]), .Y(or1res_vc_buffer31) );
    OR4X1 U2365 ( .IN1(flit31[25]), .IN2(flit31[24]), .IN3(flit31[23]), .IN4(flit31[22]), .Y(or2res_vc_buffer31) );
    OR2X1 U2366 ( .A(or1res_vc_buffer31), .B(or2res_vc_buffer31), .Y(orres_vc_buffer31) );
    AND3X1 U2367 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(norres_vc_buffer31_vc_buffer1), .IN3(orres_vc_buffer31), .Q(finres1_vc_buffer31) );
    MUX21X1 U2368 (.IN1(next_locked_vc_buffer31), .IN2(1'b1), .S(finres1_vc_buffer31), .Q(next_locked_vc_buffer31);
    AND3X1 U2369 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(flit31[33]), .IN3(flit31[32]), .Q(andres1_vc_buffer31) );
    MUX21X1 U2370 (.IN1(next_locked_vc_buffer31), .IN2(1'b0), .S(andres1_vc_buffer31), .Q(next_locked_vc_buffer31);

    INVX1 U2371 ( .A(full_vc_buffer31), .Y(full_vc_buffer31_not1) );
    INVX1 U2372 ( .A(locked_by_route_ff_vc_buffer31), .Y(locked_by_route_ff_vc_buffer31_not1) );

    MUX21X1 U2373 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer31_not1), .S(norres_vc_buffer31_vc_buffer1), .Q(thirdand_vc_buffer31);
    AND3X1 U2374 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[37]), .IN2(full_vc_buffer31_not1), .IN3(thirdand_vc_buffer31), .Q(write_flit31_vc_buffer13) );
    AND2X1 U2375 ( .IN1(full_vc_buffer31_not1), .IN2(norres_vc_buffer31_vc_buffer1), .Q(from_input_resp_input_datapath3[1]) );
    INVX1 U2376 ( .A(empty_vc_buffer31), .Y(to_output_req_in_jump_input_datapath3put_datapath3[37]) );
    AND2X1 U2377 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[37]), .IN2(to_output_resp_input_datapath3[1]), .Q(read_flit31_vc_buffer13) );
	BUFX1 U2378(.A(to_output_req_in_jump_input_datapath3put_datapath3[39:38]), .Y(2'b01));

	DFFX2 U2379 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U2380 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U2381 (.IN1(next_locked_vc_buffer31), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer31);


	BUFX1 U2382 ( .A(read_ptr_ff_fifomodule32[0]), .Y(next_read_ptr_fifomodule32[0]) );
	BUFX1 U2383 ( .A(read_ptr_ff_fifomodule32[1]), .Y(next_read_ptr_fifomodule32[1]) );
	BUFX1 U2384 ( .A(write_ptr_ff_fifomodule32[0]), .Y(next_write_ptr_fifomodule32[0]) );
	BUFX1 U2385 ( .A(write_ptr_ff_fifomodule32[1]), .Y(next_write_ptr_fifomodule32[1]) );

	XNOR2X1 U2386 ( .IN1(write_ptr_ff_fifomodule32[0]), .IN2(read_ptr_ff_fifomodule32[0]), .Q(u1temp_fifomodule32) );
	XNOR2X1 U2387 ( .IN1(write_ptr_ff_fifomodule32[1]), .IN2(read_ptr_ff_fifomodule32[1]), .Q(u2temp_fifomodule32) );
	AND2X1 U2388 ( .A(u1temp_fifomodule32), .B(u2temp_fifomodule32), .Y(empty_vc_buffer32) );
	XOR2X1 U2389 ( .A(write_ptr_ff_fifomodule32[1]), .B(read_ptr_ff_fifomodule32[1]), .Y(u4temp_fifomodule32) );
	AND2X1 U2390 ( .A(u1temp_fifomodule32), .B(u4temp_fifomodule32), .Y(full_vc_buffer32) );
	MUX21X1 U2391 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][0]));
	MUX21X1 U2392 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][1]));
	MUX21X1 U2393 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][2]));
	MUX21X1 U2394 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][3]));
	MUX21X1 U2395 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][4]));
	MUX21X1 U2396 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][5]));
	MUX21X1 U2397 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][6]));
	MUX21X1 U2398 (.IN1(fifo_ff_fifomodule32[read_ptr_ff_fifomodule32[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer32), .Q(to_output_req_in_jump_input_datapath3put_datapath3[110:77][7]));

	INVX1 U2399 ( .A(full_vc_buffer32), .Y(full_vc_buffer32_not2_fifomodule2) );
	AND2X1 U2400 ( .A(write_flit32_vc_buffer23), .B(full_vc_buffer32_not2_fifomodule2), .Y(u7temp_fifomodule32) );
	MUX21X1 U2401 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule32), .Q(u9temp_fifomodule32));
	HADDX1 U2402 ( .A0(write_ptr_ff_fifomodule32[0]), .B0(u9temp_fifomodule32), .C1(u10carry_fifomodule32), .SO(next_write_ptr_fifomodule32[0]) );
	HADDX1 U2403 ( .A0(u10carry_fifomodule32), .B0(write_ptr_ff_fifomodule32[1]), .C1(u11carry_fifomodule32), .SO(next_write_ptr_fifomodule32[1]) );

	INVX1 U2404 ( .A(empty_vc_buffer32), .Y(empty_vc_buffer32_not_fifomodule2) );
	AND2X1 U2405 ( .A(read_flit32_vc_buffer23), .B(empty_vc_buffer32_not_fifomodule2), .Y(u13temp_fifomodule32) );
	MUX21X1 U2406 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule32), .Q(u14temp_fifomodule32));
	HADDX1 U2407 ( .A0(read_ptr_ff_fifomodule32[0]), .B0(u14temp_fifomodule32), .C1(u15carry_fifomodule32), .SO(next_read_ptr_fifomodule32[0]) );
	HADDX1 U2408 ( .A0(u15carry_fifomodule32), .B0(read_ptr_ff_fifomodule32[1]), .C1(u16carry_fifomodule32), .SO(next_read_ptr_fifomodule32[1]) );

	AND2X1 U2409 ( .A(write_flit32_vc_buffer23), .B(full_vc_buffer32), .Y(u17res_fifomodule32) );
	AND2X1 U2410 ( .A(read_flit32_vc_buffer23), .B(empty_vc_buffer32), .Y(u18res_fifomodule32) );
    OR2X1 U2411 ( .A(u17res_fifomodule32), .B(u18res_fifomodule32), .Y(error_vc_buffer32) );
	XOR2X1 U2412 ( .A(write_ptr_ff_fifomodule32[0]), .B(read_ptr_ff_fifomodule32[0]), .Y(fifo_ocup_fifomodule32[0]) );
	INVX1 U2413 ( .A(write_ptr_ff_fifomodule32[0]), .Y(write_ptr_ff_fifomodule32_0_not23) );
	AND2X1 U2414 ( .A(write_ptr_ff_fifomodule32_0_not23), .B(read_ptr_ff_fifomodule32[0]), .Y(b0wire_fifomodule32) );
	XOR2X1 U2415 ( .A(write_ptr_ff_fifomodule32[1]), .B(read_ptr_ff_fifomodule32[1]), .Y(u23temp_fifomodule32) );
	INVX1 U2416 ( .A(write_ptr_ff_fifomodule32[1]), .Y(write_ptr_ff_fifomodule32_1_not23) );
	AND2X1 U2417 ( .A(read_ptr_ff_fifomodule32[1]), .B(write_ptr_ff_fifomodule32_1_not23), .Y(boutb_fifomodule32) );
	XOR2X1 U2418 ( .A(u23temp_fifomodule32), .B(b0wire_fifomodule32), .Y(fifo_ocup_fifomodule32[1]) );
	INVX1 U2419 ( .A(u23temp_fifomodule32), .Y(u23temp_fifomodule32_not_fifomodule2) );
	AND2X1 U2420 ( .A(b0wire_fifomodule32), .B(u23temp_fifomodule32_not_fifomodule2), .Y(bouta_fifomodule32) );
	OR2X1 U2421 ( .A(bouta_fifomodule32), .B(boutb_fifomodule32), .Y(boutmain_fifomodule32) );
	DFFX2 U2422 ( .CLK(clk), .D(fifo_ocup_fifomodule32[0]), .Q(ocup_o[0]) );
	DFFX2 U2423 ( .CLK(clk), .D(fifo_ocup_fifomodule32[1]), .Q(ocup_o[1]) );
	DFFX2 U2424 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule32) );
	DFFX2 U2425 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule32) );
	DFFX2 U2426 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(write_ptr_ff_fifomodule32[0]) );
	DFFX2 U2427 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(read_ptr_ff_fifomodule32[0]) );
	DFFX2 U2428 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(fifo_ff_fifomodule32[0]) );
	DFFX2 U2429 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(write_ptr_ff_fifomodule32[1]) );
	DFFX2 U2430 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(read_ptr_ff_fifomodule32[1]) );
	DFFX2 U2431 ( .CLK(arst_value_fifomodule32), .D(1'b0), .Q(fifo_ff_fifomodule32[1]) );

	DFFX2 U2432 ( .CLK(clk), .D(next_write_ptr_fifomodule32[0]), .Q(write_ptr_ff_fifomodule32[0]) );
	DFFX2 U2433 ( .CLK(clk), .D(next_write_ptr_fifomodule32[1]), .Q(write_ptr_ff_fifomodule32[1]) );
	DFFX2 U2434 ( .CLK(clk), .D(next_read_ptr_fifomodule32[0]), .Q(read_ptr_ff_fifomodule32[0]) );
	DFFX2 U2435 ( .CLK(clk), .D(next_read_ptr_fifomodule32[1]), .Q(read_ptr_ff_fifomodule32[1]) );
	  

	DFFX2 U2436 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][0]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8]) );
	DFFX2 U2437 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][1]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+1]) );
	DFFX2 U2438 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][2]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+2]) );
	DFFX2 U2439 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][3]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+3]) );
	DFFX2 U2440 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][4]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+4]) );
	DFFX2 U2441 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][5]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+5]) );
	DFFX2 U2442 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][6]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+6]) );
	DFFX2 U2443 ( .CLK(u7temp_fifomodule32), .D(from_input_req_in_jump_input_datapath3put_datapath3[110:77][7]), .Q(fifo_ff_fifomodule32[write_ptr_ff_fifomodule32[0]*8+7]) );

    BUFX1 U2444 ( .A(locked_by_route_ff_vc_buffer32), .Y(next_locked_vc_buffer32) );
    BUFX1 U2445(.A(flit32[0]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][0]));
	BUFX1 U2446(.A(flit32[1]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][1]));
	BUFX1 U2447(.A(flit32[2]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][2]));
	BUFX1 U2448(.A(flit32[3]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][3]));
	BUFX1 U2449(.A(flit32[4]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][4]));
	BUFX1 U2450(.A(flit32[5]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][5]));
	BUFX1 U2451(.A(flit32[6]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][6]));
	BUFX1 U2452(.A(flit32[7]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][7]));
	BUFX1 U2453(.A(flit32[8]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][8]));
	BUFX1 U2454(.A(flit32[9]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][9]));
	BUFX1 U2455(.A(flit32[10]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][10]));
	BUFX1 U2456(.A(flit32[11]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][11]));
	BUFX1 U2457(.A(flit32[12]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][12]));
	BUFX1 U2458(.A(flit32[13]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][13]));
	BUFX1 U2459(.A(flit32[14]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][14]));
	BUFX1 U2460(.A(flit32[15]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][15]));
	BUFX1 U2461(.A(flit32[16]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][16]));
	BUFX1 U2462(.A(flit32[17]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][17]));
	BUFX1 U2463(.A(flit32[18]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][18]));
	BUFX1 U2464(.A(flit32[19]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][19]));
	BUFX1 U2465(.A(flit32[20]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][20]));
	BUFX1 U2466(.A(flit32[21]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][21]));
	BUFX1 U2467(.A(flit32[22]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][22]));
	BUFX1 U2468(.A(flit32[23]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][23]));
	BUFX1 U2469(.A(flit32[24]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][24]));
	BUFX1 U2470(.A(flit32[25]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][25]));
	BUFX1 U2471(.A(flit32[26]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][26]));
	BUFX1 U2472(.A(flit32[27]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][27]));
	BUFX1 U2473(.A(flit32[28]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][28]));
	BUFX1 U2474(.A(flit32[29]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][29]));
	BUFX1 U2475(.A(flit32[30]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][30]));
	BUFX1 U2476(.A(flit32[31]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][31]));
	BUFX1 U2477(.A(flit32[32]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][32]));
	BUFX1 U2478(.A(flit32[33]), .Y(from_input_req_in_jump_input_datapath3put_datapath3[110:77][33]));
    NOR2X1 U2479 ( .IN1(flit32[33]), .IN2(flit32[32]), .QN(norres_vc_buffer32_vc_buffer2) );
    OR4X1 U2480 ( .IN1(flit32[29]), .IN2(flit32[28]), .IN3(flit32[27]), .IN4(flit32[26]), .Y(or1res_vc_buffer32) );
    OR4X1 U2481 ( .IN1(flit32[25]), .IN2(flit32[24]), .IN3(flit32[23]), .IN4(flit32[22]), .Y(or2res_vc_buffer32) );
    OR2X1 U2482 ( .A(or1res_vc_buffer32), .B(or2res_vc_buffer32), .Y(orres_vc_buffer32) );
    AND3X1 U2483 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(norres_vc_buffer32_vc_buffer2), .IN3(orres_vc_buffer32), .Q(finres1_vc_buffer32) );
    MUX21X1 U2484 (.IN1(next_locked_vc_buffer32), .IN2(1'b1), .S(finres1_vc_buffer32), .Q(next_locked_vc_buffer32);
    AND3X1 U2485 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(flit32[33]), .IN3(flit32[32]), .Q(andres1_vc_buffer32) );
    MUX21X1 U2486 (.IN1(next_locked_vc_buffer32), .IN2(1'b0), .S(andres1_vc_buffer32), .Q(next_locked_vc_buffer32);

    INVX1 U2487 ( .A(full_vc_buffer32), .Y(full_vc_buffer32_not2) );
    INVX1 U2488 ( .A(locked_by_route_ff_vc_buffer32), .Y(locked_by_route_ff_vc_buffer32_not2) );

    MUX21X1 U2489 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer32_not2), .S(norres_vc_buffer32_vc_buffer2), .Q(thirdand_vc_buffer32);
    AND3X1 U2490 ( .IN1(from_input_req_in_jump_input_datapath3put_datapath3[74]), .IN2(full_vc_buffer32_not2), .IN3(thirdand_vc_buffer32), .Q(write_flit32_vc_buffer23) );
    AND2X1 U2491 ( .IN1(full_vc_buffer32_not2), .IN2(norres_vc_buffer32_vc_buffer2), .Q(from_input_resp_input_datapath3[2]) );
    INVX1 U2492 ( .A(empty_vc_buffer32), .Y(to_output_req_in_jump_input_datapath3put_datapath3[74]) );
    AND2X1 U2493 ( .IN1(to_output_req_in_jump_input_datapath3put_datapath3[74]), .IN2(to_output_resp_input_datapath3[2]), .Q(read_flit32_vc_buffer23) );
	BUFX1 U2494(.A(to_output_req_in_jump_input_datapath3put_datapath3[76:75]), .Y(2'b10));

	DFFX2 U2495 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U2496 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U2497 (.IN1(next_locked_vc_buffer32), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer32);

	BUFX1 U2498(.A(from_input_req_in_jump_input_datapath3put_datapath3[77]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U2499(.A(from_input_req_in_jump_input_datapath3put_datapath3[78]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U2500(.A(from_input_req_in_jump_input_datapath3put_datapath3[79]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U2501(.A(from_input_req_in_jump_input_datapath3put_datapath3[80]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U2502(.A(from_input_req_in_jump_input_datapath3put_datapath3[81]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U2503(.A(from_input_req_in_jump_input_datapath3put_datapath3[82]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U2504(.A(from_input_req_in_jump_input_datapath3put_datapath3[83]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U2505(.A(from_input_req_in_jump_input_datapath3put_datapath3[84]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U2506(.A(from_input_req_in_jump_input_datapath3put_datapath3[85]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U2507(.A(from_input_req_in_jump_input_datapath3put_datapath3[86]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U2508(.A(from_input_req_in_jump_input_datapath3put_datapath3[87]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U2509(.A(from_input_req_in_jump_input_datapath3put_datapath3[88]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U2510(.A(from_input_req_in_jump_input_datapath3put_datapath3[89]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U2511(.A(from_input_req_in_jump_input_datapath3put_datapath3[90]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U2512(.A(from_input_req_in_jump_input_datapath3put_datapath3[91]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U2513(.A(from_input_req_in_jump_input_datapath3put_datapath3[92]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U2514(.A(from_input_req_in_jump_input_datapath3put_datapath3[93]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U2515(.A(from_input_req_in_jump_input_datapath3put_datapath3[94]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U2516(.A(from_input_req_in_jump_input_datapath3put_datapath3[95]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U2517(.A(from_input_req_in_jump_input_datapath3put_datapath3[96]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U2518(.A(from_input_req_in_jump_input_datapath3put_datapath3[97]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U2519(.A(from_input_req_in_jump_input_datapath3put_datapath3[98]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U2520(.A(from_input_req_in_jump_input_datapath3put_datapath3[99]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U2521(.A(from_input_req_in_jump_input_datapath3put_datapath3[100]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U2522(.A(from_input_req_in_jump_input_datapath3put_datapath3[101]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U2523(.A(from_input_req_in_jump_input_datapath3put_datapath3[102]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U2524(.A(from_input_req_in_jump_input_datapath3put_datapath3[103]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U2525(.A(from_input_req_in_jump_input_datapath3put_datapath3[104]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U2526(.A(from_input_req_in_jump_input_datapath3put_datapath3[105]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U2527(.A(from_input_req_in_jump_input_datapath3put_datapath3[106]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U2528(.A(from_input_req_in_jump_input_datapath3put_datapath3[107]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U2529(.A(from_input_req_in_jump_input_datapath3put_datapath3[108]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U2530(.A(from_input_req_in_jump_input_datapath3put_datapath3[109]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U2531(.A(from_input_req_in_jump_input_datapath3put_datapath3[110]), .Y(ext_req_v_i[147:111][36]));
    XNOR2X1 U2532 ( .IN1(ext_req_v_i[147:111][1]), .IN2(i_input_datapath3[0]), .QN(xnor1resu_input_datapath3) );
    XNOR2X1 U2533 ( .IN1(ext_req_v_i[147:111][2]), .IN2(i_input_datapath3[1]), .QN(xnor2resu_input_datapath3) );
    AND2X1 U2534 ( .IN1(xnor1resu_input_datapath3), .IN2(xnor2resu_input_datapath3), .Q(and1resu_input_datapath3) );
    AND3X1 U2535 ( .IN1(and1resu_input_datapath3), .IN2(ext_req_v_i[147:111][0]), .IN2(ext_req_v_i[147:111][0]), .Q(cond1line_input_datapath3) );
    MUX21X1 U2536 (.IN1(vc_ch_act_in_input_datapath3[0]), .IN2(i_input_datapath3[0]), .S(cond1line_input_datapath3), .Q(vc_ch_act_in_input_datapath3[0]));
    MUX21X1 U2537 (.IN1(vc_ch_act_in_input_datapath3[1]), .IN2(i_input_datapath3[1]), .S(cond1line_input_datapath3), .Q(vc_ch_act_in_input_datapath3[1]));
    MUX21X1 U2538 (.IN1(req_in_jump_input_datapath3), .IN2(1), .S(cond1line_input_datapath3), .Q(req_in_jump_input_datapath3));
	BUFX1 U2539(.A(from_input_req_in_jump_input_datapath3put_datapath3[40]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U2540(.A(from_input_req_in_jump_input_datapath3put_datapath3[41]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U2541(.A(from_input_req_in_jump_input_datapath3put_datapath3[42]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U2542(.A(from_input_req_in_jump_input_datapath3put_datapath3[43]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U2543(.A(from_input_req_in_jump_input_datapath3put_datapath3[44]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U2544(.A(from_input_req_in_jump_input_datapath3put_datapath3[45]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U2545(.A(from_input_req_in_jump_input_datapath3put_datapath3[46]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U2546(.A(from_input_req_in_jump_input_datapath3put_datapath3[47]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U2547(.A(from_input_req_in_jump_input_datapath3put_datapath3[48]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U2548(.A(from_input_req_in_jump_input_datapath3put_datapath3[49]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U2549(.A(from_input_req_in_jump_input_datapath3put_datapath3[50]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U2550(.A(from_input_req_in_jump_input_datapath3put_datapath3[51]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U2551(.A(from_input_req_in_jump_input_datapath3put_datapath3[52]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U2552(.A(from_input_req_in_jump_input_datapath3put_datapath3[53]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U2553(.A(from_input_req_in_jump_input_datapath3put_datapath3[54]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U2554(.A(from_input_req_in_jump_input_datapath3put_datapath3[55]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U2555(.A(from_input_req_in_jump_input_datapath3put_datapath3[56]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U2556(.A(from_input_req_in_jump_input_datapath3put_datapath3[57]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U2557(.A(from_input_req_in_jump_input_datapath3put_datapath3[58]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U2558(.A(from_input_req_in_jump_input_datapath3put_datapath3[59]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U2559(.A(from_input_req_in_jump_input_datapath3put_datapath3[60]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U2560(.A(from_input_req_in_jump_input_datapath3put_datapath3[61]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U2561(.A(from_input_req_in_jump_input_datapath3put_datapath3[62]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U2562(.A(from_input_req_in_jump_input_datapath3put_datapath3[63]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U2563(.A(from_input_req_in_jump_input_datapath3put_datapath3[64]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U2564(.A(from_input_req_in_jump_input_datapath3put_datapath3[65]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U2565(.A(from_input_req_in_jump_input_datapath3put_datapath3[66]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U2566(.A(from_input_req_in_jump_input_datapath3put_datapath3[67]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U2567(.A(from_input_req_in_jump_input_datapath3put_datapath3[68]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U2568(.A(from_input_req_in_jump_input_datapath3put_datapath3[69]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U2569(.A(from_input_req_in_jump_input_datapath3put_datapath3[70]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U2570(.A(from_input_req_in_jump_input_datapath3put_datapath3[71]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U2571(.A(from_input_req_in_jump_input_datapath3put_datapath3[72]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U2572(.A(from_input_req_in_jump_input_datapath3put_datapath3[73]), .Y(ext_req_v_i[147:111][36]));

	BUFX1 U2573(.A(from_input_req_in_jump_input_datapath3put_datapath3[3]), .Y(ext_req_v_i[147:111][3]));
	BUFX1 U2574(.A(from_input_req_in_jump_input_datapath3put_datapath3[4]), .Y(ext_req_v_i[147:111][4]));
	BUFX1 U2575(.A(from_input_req_in_jump_input_datapath3put_datapath3[5]), .Y(ext_req_v_i[147:111][5]));
	BUFX1 U2576(.A(from_input_req_in_jump_input_datapath3put_datapath3[6]), .Y(ext_req_v_i[147:111][6]));
	BUFX1 U2577(.A(from_input_req_in_jump_input_datapath3put_datapath3[7]), .Y(ext_req_v_i[147:111][7]));
	BUFX1 U2578(.A(from_input_req_in_jump_input_datapath3put_datapath3[8]), .Y(ext_req_v_i[147:111][8]));
	BUFX1 U2579(.A(from_input_req_in_jump_input_datapath3put_datapath3[9]), .Y(ext_req_v_i[147:111][9]));
	BUFX1 U2580(.A(from_input_req_in_jump_input_datapath3put_datapath3[10]), .Y(ext_req_v_i[147:111][10]));
	BUFX1 U2581(.A(from_input_req_in_jump_input_datapath3put_datapath3[11]), .Y(ext_req_v_i[147:111][11]));
	BUFX1 U2582(.A(from_input_req_in_jump_input_datapath3put_datapath3[12]), .Y(ext_req_v_i[147:111][12]));
	BUFX1 U2583(.A(from_input_req_in_jump_input_datapath3put_datapath3[13]), .Y(ext_req_v_i[147:111][13]));
	BUFX1 U2584(.A(from_input_req_in_jump_input_datapath3put_datapath3[14]), .Y(ext_req_v_i[147:111][14]));
	BUFX1 U2585(.A(from_input_req_in_jump_input_datapath3put_datapath3[15]), .Y(ext_req_v_i[147:111][15]));
	BUFX1 U2586(.A(from_input_req_in_jump_input_datapath3put_datapath3[16]), .Y(ext_req_v_i[147:111][16]));
	BUFX1 U2587(.A(from_input_req_in_jump_input_datapath3put_datapath3[17]), .Y(ext_req_v_i[147:111][17]));
	BUFX1 U2588(.A(from_input_req_in_jump_input_datapath3put_datapath3[18]), .Y(ext_req_v_i[147:111][18]));
	BUFX1 U2589(.A(from_input_req_in_jump_input_datapath3put_datapath3[19]), .Y(ext_req_v_i[147:111][19]));
	BUFX1 U2590(.A(from_input_req_in_jump_input_datapath3put_datapath3[20]), .Y(ext_req_v_i[147:111][20]));
	BUFX1 U2591(.A(from_input_req_in_jump_input_datapath3put_datapath3[21]), .Y(ext_req_v_i[147:111][21]));
	BUFX1 U2592(.A(from_input_req_in_jump_input_datapath3put_datapath3[22]), .Y(ext_req_v_i[147:111][22]));
	BUFX1 U2593(.A(from_input_req_in_jump_input_datapath3put_datapath3[23]), .Y(ext_req_v_i[147:111][23]));
	BUFX1 U2594(.A(from_input_req_in_jump_input_datapath3put_datapath3[24]), .Y(ext_req_v_i[147:111][24]));
	BUFX1 U2595(.A(from_input_req_in_jump_input_datapath3put_datapath3[25]), .Y(ext_req_v_i[147:111][25]));
	BUFX1 U2596(.A(from_input_req_in_jump_input_datapath3put_datapath3[26]), .Y(ext_req_v_i[147:111][26]));
	BUFX1 U2597(.A(from_input_req_in_jump_input_datapath3put_datapath3[27]), .Y(ext_req_v_i[147:111][27]));
	BUFX1 U2598(.A(from_input_req_in_jump_input_datapath3put_datapath3[28]), .Y(ext_req_v_i[147:111][28]));
	BUFX1 U2599(.A(from_input_req_in_jump_input_datapath3put_datapath3[29]), .Y(ext_req_v_i[147:111][29]));
	BUFX1 U2600(.A(from_input_req_in_jump_input_datapath3put_datapath3[30]), .Y(ext_req_v_i[147:111][30]));
	BUFX1 U2601(.A(from_input_req_in_jump_input_datapath3put_datapath3[31]), .Y(ext_req_v_i[147:111][31]));
	BUFX1 U2602(.A(from_input_req_in_jump_input_datapath3put_datapath3[32]), .Y(ext_req_v_i[147:111][32]));
	BUFX1 U2603(.A(from_input_req_in_jump_input_datapath3put_datapath3[33]), .Y(ext_req_v_i[147:111][33]));
	BUFX1 U2604(.A(from_input_req_in_jump_input_datapath3put_datapath3[34]), .Y(ext_req_v_i[147:111][34]));
	BUFX1 U2605(.A(from_input_req_in_jump_input_datapath3put_datapath3[35]), .Y(ext_req_v_i[147:111][35]));
	BUFX1 U2606(.A(from_input_req_in_jump_input_datapath3put_datapath3[36]), .Y(ext_req_v_i[147:111][36]));

    MUX21X1 U2607 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3 * 37]), .IN2(ext_req_v_i[147:111][0]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3 * 37]));
    MUX21X1 U2608 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+2]), .IN2(vc_ch_act_in_input_datapath3[1]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+2]));
    MUX21X1 U2609 (.IN1(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+1]), .IN2(vc_ch_act_in_input_datapath3[0]), .S(req_in_jump_input_datapath3), .Q(from_input_req_in_jump_input_datapath3put_datapath3[vc_ch_act_in_input_datapath3*37+1]));
    MUX21X1 U2610 (.IN1(ext_resp_v_o[4:3][0]), .IN2(from_input_resp_input_datapath3[vc_ch_act_in_input_datapath3]), .S(req_in_jump_input_datapath3), .Q(ext_resp_v_o[4:3][0]));

    INVX1 U2611 ( .A(req_in_jump_input_datapath3), .Y(req_in_jump_input_datapath3_not) );
    MUX21X1 U2612 (.IN1(ext_resp_v_o[4:3][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath3_not), .Q(ext_resp_v_o[4:3][0]));
    BUFX1 U2613(.A(from_input_req_in_jump_input_datapath3put_datapath3[34]), .Y(ext_req_v_i[147:111][34]));

    XOR2X1 U2614 ( .IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b1), .Q(xor1resu_input_datapath3) );
    MUX21X1 U2615 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(xor1resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U2616 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b0), .S(xor1resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[1]));
    AND2X1 U2617 ( .IN1(xor1resu_input_datapath3), .IN2(to_output_req_in_jump_input_datapath3put_datapath3[j_input_datapath3*37]), .Q(and2resu_input_datapath3) );
    MUX21X1 U2618 (.IN1(vc_ch_act_out_input_datapath3[0]), .IN2(j_input_datapath3[0]), .S(and2resu_input_datapath3), .Q(vc_ch_act_out_input_datapath3[0]));
    MUX21X1 U2619 (.IN1(vc_ch_act_out_input_datapath3[1]), .IN2(j_input_datapath3[1]), .S(and2resu_input_datapath3), .Q(vc_ch_act_out_input_datapath3[1]));
    MUX21X1 U2620 (.IN1(req_out_jump_input_datapath3), .IN2(1'b1), .S(and2resu_input_datapath3), .Q(req_out_jump_input_datapath3));
    MUX21X1 U2621 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(and2resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U2622 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b1), .S(and2resu_input_datapath3), .Q(_sv2v_jump_input_datapath3[1]));
    HADDX1 U2623 ( .A0(j_input_datapath3[0]), .B0(1'b1), .C1(j_input_datapath3[1]), .SO(j_input_datapath3[0]) );
    HADDX1 U2624 ( .A0(j_input_datapath3[0]), .B0(1'b1), .C1(j_input_datapath3[1]), .SO(j_input_datapath3[0]) );
    AND2X1 U2625 ( .IN1(xor1resu_input_datapath3), .IN2(to_output_req_in_jump_input_datapath3put_datapath3[j_input_datapath3*37]), .Q(and3resu) );
    NAND2X1 U2626(.A(_sv2v_jump_input_datapath3[0]),.B(_sv2v_jump_input_datapath3[1]),.Y(nand1resu_input_datapath33));
    MUX21X1 U2627 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(1'b0), .S(nand1resu_input_datapath33), .Q(_sv2v_jump_input_datapath3[0]));
    MUX21X1 U2628 (.IN1(_sv2v_jump_input_datapath3[1]), .IN2(1'b0), .S(nand1resu_input_datapath33), .Q(_sv2v_jump_input_datapath3[1]));
    XNOR2X1 U2629 (.IN1(_sv2v_jump_input_datapath3[0]), .IN2(_sv2v_jump_input_datapath3[1]), .Q(xnor23resu_input_datapath3) );
    AND2X1 U2630 ( .IN1(xnor23resu_input_datapath3), .IN2(req_out_jump_input_datapath3), .Q(and4resu_input_datapath3) );

    MUX21X1 U2631(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[147:111][3]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U2632(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[147:111][4]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U2633(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[147:111][5]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U2634(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[147:111][6]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U2635(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[147:111][7]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U2636(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[147:111][8]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U2637(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[147:111][9]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U2638(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[147:111][10]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U2639(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[147:111][11]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U2640(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[147:111][12]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U2641(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[147:111][13]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U2642(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[147:111][14]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U2643(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[147:111][15]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U2644(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[147:111][16]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U2645(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[147:111][17]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U2646(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[147:111][18]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U2647(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[147:111][19]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U2648(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[147:111][20]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U2649(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[147:111][21]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U2650(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[147:111][22]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U2651(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[147:111][23]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U2652(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[147:111][24]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U2653(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[147:111][25]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U2654(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[147:111][26]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U2655(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[147:111][27]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U2656(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[147:111][28]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U2657(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[147:111][29]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U2658(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[147:111][30]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U2659(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[147:111][31]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U2660(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[147:111][32]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U2661(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[147:111][33]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U2662(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[147:111][34]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U2663(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[147:111][35]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U2664(.IN1(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[147:111][36]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U2665(.IN1(int_req_v[147:111][0]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3 * 37)]), .S(and4resu_input_datapath3), .Q(int_req_v[147:111][0]));
	MUX21X1 U2666(.IN1(int_req_v[147:111][1]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+1]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+1]));
	MUX21X1 U2667(.IN1(int_req_v[147:111][2]),.IN2(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+2]), .S(and4resu_input_datapath3), .Q(to_output_req_in_jump_input_datapath3put_datapath3[(vc_ch_act_out_input_datapath3*37)+2]));
	MUX21X1 U2668(.IN1(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3]),.IN2(int_resp_v[4:3]), .S(and4resu_input_datapath3), .Q(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3]));
	MUX21X1 U2669(.IN1(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3+1]),.IN2(int_resp_v[4:3]), .S(and4resu_input_datapath3), .Q(to_output_resp_input_datapath3[vc_ch_act_out_input_datapath3+1]));

	BUFX1 U2670 ( .A(read_ptr_ff_fifomodule4[0]), .Y(next_read_ptr_fifomodule4[0]) );
	BUFX1 U2671 ( .A(read_ptr_ff_fifomodule4[1]), .Y(next_read_ptr_fifomodule4[1]) );
	BUFX1 U2672 ( .A(write_ptr_ff_fifomodule4[0]), .Y(next_write_ptr_fifomodule4[0]) );
	BUFX1 U2673 ( .A(write_ptr_ff_fifomodule4[1]), .Y(next_write_ptr_fifomodule4[1]) );

	XNOR2X1 U2674 ( .IN1(write_ptr_ff_fifomodule4[0]), .IN2(read_ptr_ff_fifomodule4[0]), .Q(u1temp_fifomodule4) );
	XNOR2X1 U2675 ( .IN1(write_ptr_ff_fifomodule4[1]), .IN2(read_ptr_ff_fifomodule4[1]), .Q(u2temp_fifomodule4) );
	AND2X1 U2676 ( .A(u1temp_fifomodule4), .B(u2temp_fifomodule4), .Y(empty_vc_buffer4) );
	XOR2X1 U2677 ( .A(write_ptr_ff_fifomodule4[1]), .B(read_ptr_ff_fifomodule4[1]), .Y(u4temp_fifomodule4) );
	AND2X1 U2678 ( .A(u1temp_fifomodule4), .B(u4temp_fifomodule4), .Y(full_vc_buffer4) );
	MUX21X1 U2679 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][0]));
	MUX21X1 U2680 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][1]));
	MUX21X1 U2681 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][2]));
	MUX21X1 U2682 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][3]));
	MUX21X1 U2683 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][4]));
	MUX21X1 U2684 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][5]));
	MUX21X1 U2685 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][6]));
	MUX21X1 U2686 (.IN1(fifo_ff_fifomodule4[read_ptr_ff_fifomodule4[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[36:3][7]));

	INVX1 U2687 ( .A(full_vc_buffer4), .Y(full_vc_buffer4_not_fifomodule) );
	AND2X1 U2688 ( .A(write_flit4_vc_buffer4), .B(full_vc_buffer4_not_fifomodule), .Y(u7temp_fifomodule4) );
	MUX21X1 U2689 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule4), .Q(u9temp_fifomodule4));
	HADDX1 U2690 ( .A0(write_ptr_ff_fifomodule4[0]), .B0(u9temp_fifomodule4), .C1(u10carry_fifomodule4), .SO(next_write_ptr_fifomodule4[0]) );
	HADDX1 U2691 ( .A0(u10carry_fifomodule4), .B0(write_ptr_ff_fifomodule4[1]), .C1(u11carry_fifomodule4), .SO(next_write_ptr_fifomodule4[1]) );

	INVX1 U2692 ( .A(empty_vc_buffer4), .Y(empty_vc_buffer4_not_fifomodule) );
	AND2X1 U2693 ( .A(read_flit4_vc_buffer4), .B(empty_vc_buffer4_not_fifomodule), .Y(u13temp_fifomodule4) );
	MUX21X1 U2694 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule4), .Q(u14temp_fifomodule4));
	HADDX1 U2695 ( .A0(read_ptr_ff_fifomodule4[0]), .B0(u14temp_fifomodule4), .C1(u15carry_fifomodule4), .SO(next_read_ptr_fifomodule4[0]) );
	HADDX1 U2696 ( .A0(u15carry_fifomodule4), .B0(read_ptr_ff_fifomodule4[1]), .C1(u16carry_fifomodule4), .SO(next_read_ptr_fifomodule4[1]) );

	AND2X1 U2697 ( .A(write_flit4_vc_buffer4), .B(full_vc_buffer4), .Y(u17res_fifomodule4) );
	AND2X1 U2698 ( .A(read_flit4_vc_buffer4), .B(empty_vc_buffer4), .Y(u18res_fifomodule4) );
    OR2X1 U2699 ( .A(u17res_fifomodule4), .B(u18res_fifomodule4), .Y(error_vc_buffer4) );
	XOR2X1 U2700 ( .A(write_ptr_ff_fifomodule4[0]), .B(read_ptr_ff_fifomodule4[0]), .Y(fifo_ocup_fifomodule4[0]) );
	INVX1 U2701 ( .A(write_ptr_ff_fifomodule4[0]), .Y(write_ptr_ff_fifomodule4_0_not4) );
	AND2X1 U2702 ( .A(write_ptr_ff_fifomodule4_0_not4), .B(read_ptr_ff_fifomodule4[0]), .Y(b0wire_fifomodule4) );
	XOR2X1 U2703 ( .A(write_ptr_ff_fifomodule4[1]), .B(read_ptr_ff_fifomodule4[1]), .Y(u23temp_fifomodule4) );
	INVX1 U2704 ( .A(write_ptr_ff_fifomodule4[1]), .Y(write_ptr_ff_fifomodule4_1_not4) );
	AND2X1 U2705 ( .A(read_ptr_ff_fifomodule4[1]), .B(write_ptr_ff_fifomodule4_1_not4), .Y(boutb_fifomodule4) );
	XOR2X1 U2706 ( .A(u23temp_fifomodule4), .B(b0wire_fifomodule4), .Y(fifo_ocup_fifomodule4[1]) );
	INVX1 U2707 ( .A(u23temp_fifomodule4), .Y(u23temp_fifomodule4_not_fifomodule4) );
	AND2X1 U2708 ( .A(b0wire_fifomodule4), .B(u23temp_fifomodule4_not_fifomodule4), .Y(bouta_fifomodule4) );
	OR2X1 U2709 ( .A(bouta_fifomodule4), .B(boutb_fifomodule4), .Y(boutmain_fifomodule4) );
	DFFX2 U2710 ( .CLK(clk), .D(fifo_ocup_fifomodule4[0]), .Q(ocup_o[0]) );
	DFFX2 U2711 ( .CLK(clk), .D(fifo_ocup_fifomodule4[1]), .Q(ocup_o[1]) );
	DFFX2 U2712 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule4) );
	DFFX2 U2713 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule4) );
	DFFX2 U2714 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(write_ptr_ff_fifomodule4[0]) );
	DFFX2 U2715 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(read_ptr_ff_fifomodule4[0]) );
	DFFX2 U2716 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(fifo_ff_fifomodule4[0]) );
	DFFX2 U2717 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(write_ptr_ff_fifomodule4[1]) );
	DFFX2 U2718 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(read_ptr_ff_fifomodule4[1]) );
	DFFX2 U2719 ( .CLK(arst_value_fifomodule4), .D(1'b0), .Q(fifo_ff_fifomodule4[1]) );

	DFFX2 U2720 ( .CLK(clk), .D(next_write_ptr_fifomodule4[0]), .Q(write_ptr_ff_fifomodule4[0]) );
	DFFX2 U2721 ( .CLK(clk), .D(next_write_ptr_fifomodule4[1]), .Q(write_ptr_ff_fifomodule4[1]) );
	DFFX2 U2722 ( .CLK(clk), .D(next_read_ptr_fifomodule4[0]), .Q(read_ptr_ff_fifomodule4[0]) );
	DFFX2 U2723 ( .CLK(clk), .D(next_read_ptr_fifomodule4[1]), .Q(read_ptr_ff_fifomodule4[1]) );
	  

	DFFX2 U2724 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][0]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8]) );
	DFFX2 U2725 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][1]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+1]) );
	DFFX2 U2726 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][2]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+2]) );
	DFFX2 U2727 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][3]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+3]) );
	DFFX2 U2728 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][4]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+4]) );
	DFFX2 U2729 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][5]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+5]) );
	DFFX2 U2730 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][6]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+6]) );
	DFFX2 U2731 ( .CLK(u7temp_fifomodule4), .D(from_input_req_in_jump_input_datapath4put_datapath4[36:3][7]), .Q(fifo_ff_fifomodule4[write_ptr_ff_fifomodule4[0]*8+7]) );

    BUFX1 U2732 ( .A(locked_by_route_ff_vc_buffer4), .Y(next_locked_vc_buffer4) );
    BUFX1 U2733(.A(flit4[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][0]));
	BUFX1 U2734(.A(flit4[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][1]));
	BUFX1 U2735(.A(flit4[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][2]));
	BUFX1 U2736(.A(flit4[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][3]));
	BUFX1 U2737(.A(flit4[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][4]));
	BUFX1 U2738(.A(flit4[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][5]));
	BUFX1 U2739(.A(flit4[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][6]));
	BUFX1 U2740(.A(flit4[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][7]));
	BUFX1 U2741(.A(flit4[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][8]));
	BUFX1 U2742(.A(flit4[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][9]));
	BUFX1 U2743(.A(flit4[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][10]));
	BUFX1 U2744(.A(flit4[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][11]));
	BUFX1 U2745(.A(flit4[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][12]));
	BUFX1 U2746(.A(flit4[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][13]));
	BUFX1 U2747(.A(flit4[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][14]));
	BUFX1 U2748(.A(flit4[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][15]));
	BUFX1 U2749(.A(flit4[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][16]));
	BUFX1 U2750(.A(flit4[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][17]));
	BUFX1 U2751(.A(flit4[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][18]));
	BUFX1 U2752(.A(flit4[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][19]));
	BUFX1 U2753(.A(flit4[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][20]));
	BUFX1 U2754(.A(flit4[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][21]));
	BUFX1 U2755(.A(flit4[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][22]));
	BUFX1 U2756(.A(flit4[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][23]));
	BUFX1 U2757(.A(flit4[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][24]));
	BUFX1 U2758(.A(flit4[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][25]));
	BUFX1 U2759(.A(flit4[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][26]));
	BUFX1 U2760(.A(flit4[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][27]));
	BUFX1 U2761(.A(flit4[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][28]));
	BUFX1 U2762(.A(flit4[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][29]));
	BUFX1 U2763(.A(flit4[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][30]));
	BUFX1 U2764(.A(flit4[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][31]));
	BUFX1 U2765(.A(flit4[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][32]));
	BUFX1 U2766(.A(flit4[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[36:3][33]));
    NOR2X1 U2767 ( .IN1(flit4[33]), .IN2(flit4[32]), .QN(norres_vc_buffer4_vc_buffer4) );
    OR4X1 U2768 ( .IN1(flit4[29]), .IN2(flit4[28]), .IN3(flit4[27]), .IN4(flit4[26]), .Y(or1res_vc_buffer4) );
    OR4X1 U2769 ( .IN1(flit4[25]), .IN2(flit4[24]), .IN3(flit4[23]), .IN4(flit4[22]), .Y(or2res_vc_buffer4) );
    OR2X1 U2770 ( .A(or1res_vc_buffer4), .B(or2res_vc_buffer4), .Y(orres_vc_buffer4) );
    AND3X1 U2771 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(norres_vc_buffer4_vc_buffer4), .IN3(orres_vc_buffer4), .Q(finres1_vc_buffer4) );
    MUX21X1 U2772 (.IN1(next_locked_vc_buffer4), .IN2(1'b1), .S(finres1_vc_buffer4), .Q(next_locked_vc_buffer4);
    AND3X1 U2773 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(flit4[33]), .IN3(flit4[32]), .Q(andres1_vc_buffer4) );
    MUX21X1 U2774 (.IN1(next_locked_vc_buffer4), .IN2(1'b0), .S(andres1_vc_buffer4), .Q(next_locked_vc_buffer4);

    INVX1 U2775 ( .A(full_vc_buffer4), .Y(full_vc_buffer4_not) );
    INVX1 U2776 ( .A(locked_by_route_ff_vc_buffer4), .Y(locked_by_route_ff_vc_buffer4_not) );

    MUX21X1 U2777 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer4_not), .S(norres_vc_buffer4_vc_buffer4), .Q(thirdand_vc_buffer4);
    AND3X1 U2778 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[0]), .IN2(full_vc_buffer4_not), .IN3(thirdand_vc_buffer4), .Q(write_flit4_vc_buffer4) );
    AND2X1 U2779 ( .IN1(full_vc_buffer4_not), .IN2(norres_vc_buffer4_vc_buffer4), .Q(from_input_resp_input_datapath4[0]) );
    INVX1 U2780 ( .A(empty_vc_buffer4), .Y(to_output_req_in_jump_input_datapath4put_datapath4[0]) );
    AND2X1 U2781 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[0]), .IN2(to_output_resp_input_datapath4[0]), .Q(read_flit4_vc_buffer4) );
	BUFX1 U2782(.A(to_output_req_in_jump_input_datapath4put_datapath4[2:1]), .Y(2'b00));

	DFFX2 U2783 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U2784 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U2785 (.IN1(next_locked_vc_buffer4), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer4);

	BUFX1 U2786 ( .A(read_ptr_ff_fifomodule41[0]), .Y(next_read_ptr_fifomodule41[0]) );
	BUFX1 U2787 ( .A(read_ptr_ff_fifomodule41[1]), .Y(next_read_ptr_fifomodule41[1]) );
	BUFX1 U2788 ( .A(write_ptr_ff_fifomodule41[0]), .Y(next_write_ptr_fifomodule41[0]) );
	BUFX1 U2789 ( .A(write_ptr_ff_fifomodule41[1]), .Y(next_write_ptr_fifomodule41[1]) );

	XNOR2X1 U2790 ( .IN1(write_ptr_ff_fifomodule41[0]), .IN2(read_ptr_ff_fifomodule41[0]), .Q(u1temp_fifomodule41) );
	XNOR2X1 U2791 ( .IN1(write_ptr_ff_fifomodule41[1]), .IN2(read_ptr_ff_fifomodule41[1]), .Q(u2temp_fifomodule41) );
	AND2X1 U2792 ( .A(u1temp_fifomodule41), .B(u2temp_fifomodule41), .Y(empty_vc_buffer41) );
	XOR2X1 U2793 ( .A(write_ptr_ff_fifomodule41[1]), .B(read_ptr_ff_fifomodule41[1]), .Y(u4temp_fifomodule41) );
	AND2X1 U2794 ( .A(u1temp_fifomodule41), .B(u4temp_fifomodule41), .Y(full_vc_buffer41) );
	MUX21X1 U2795 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][0]));
	MUX21X1 U2796 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][1]));
	MUX21X1 U2797 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][2]));
	MUX21X1 U2798 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][3]));
	MUX21X1 U2799 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][4]));
	MUX21X1 U2800 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][5]));
	MUX21X1 U2801 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][6]));
	MUX21X1 U2802 (.IN1(fifo_ff_fifomodule41[read_ptr_ff_fifomodule41[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer41), .Q(to_output_req_in_jump_input_datapath4put_datapath4[73:40][7]));

	INVX1 U2803 ( .A(full_vc_buffer41), .Y(full_vc_buffer41_not1_fifomodule1) );
	AND2X1 U2804 ( .A(write_flit41_vc_buffer14), .B(full_vc_buffer41_not1_fifomodule1), .Y(u7temp_fifomodule41) );
	MUX21X1 U2805 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule41), .Q(u9temp_fifomodule41));
	HADDX1 U2806 ( .A0(write_ptr_ff_fifomodule41[0]), .B0(u9temp_fifomodule41), .C1(u10carry_fifomodule41), .SO(next_write_ptr_fifomodule41[0]) );
	HADDX1 U2807 ( .A0(u10carry_fifomodule41), .B0(write_ptr_ff_fifomodule41[1]), .C1(u11carry_fifomodule41), .SO(next_write_ptr_fifomodule41[1]) );

	INVX1 U2808 ( .A(empty_vc_buffer41), .Y(empty_vc_buffer41_not_fifomodule1) );
	AND2X1 U2809 ( .A(read_flit41_vc_buffer14), .B(empty_vc_buffer41_not_fifomodule1), .Y(u13temp_fifomodule41) );
	MUX21X1 U2810 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule41), .Q(u14temp_fifomodule41));
	HADDX1 U2811 ( .A0(read_ptr_ff_fifomodule41[0]), .B0(u14temp_fifomodule41), .C1(u15carry_fifomodule41), .SO(next_read_ptr_fifomodule41[0]) );
	HADDX1 U2812 ( .A0(u15carry_fifomodule41), .B0(read_ptr_ff_fifomodule41[1]), .C1(u16carry_fifomodule41), .SO(next_read_ptr_fifomodule41[1]) );

	AND2X1 U2813 ( .A(write_flit41_vc_buffer14), .B(full_vc_buffer41), .Y(u17res_fifomodule41) );
	AND2X1 U2814 ( .A(read_flit41_vc_buffer14), .B(empty_vc_buffer41), .Y(u18res_fifomodule41) );
    OR2X1 U2815 ( .A(u17res_fifomodule41), .B(u18res_fifomodule41), .Y(error_vc_buffer41) );
	XOR2X1 U2816 ( .A(write_ptr_ff_fifomodule41[0]), .B(read_ptr_ff_fifomodule41[0]), .Y(fifo_ocup_fifomodule41[0]) );
	INVX1 U2817 ( .A(write_ptr_ff_fifomodule41[0]), .Y(write_ptr_ff_fifomodule41_0_not14) );
	AND2X1 U2818 ( .A(write_ptr_ff_fifomodule41_0_not14), .B(read_ptr_ff_fifomodule41[0]), .Y(b0wire_fifomodule41) );
	XOR2X1 U2819 ( .A(write_ptr_ff_fifomodule41[1]), .B(read_ptr_ff_fifomodule41[1]), .Y(u23temp_fifomodule41) );
	INVX1 U2820 ( .A(write_ptr_ff_fifomodule41[1]), .Y(write_ptr_ff_fifomodule41_1_not14) );
	AND2X1 U2821 ( .A(read_ptr_ff_fifomodule41[1]), .B(write_ptr_ff_fifomodule41_1_not14), .Y(boutb_fifomodule41) );
	XOR2X1 U2822 ( .A(u23temp_fifomodule41), .B(b0wire_fifomodule41), .Y(fifo_ocup_fifomodule41[1]) );
	INVX1 U2823 ( .A(u23temp_fifomodule41), .Y(u23temp_fifomodule41_not_fifomodule1) );
	AND2X1 U2824 ( .A(b0wire_fifomodule41), .B(u23temp_fifomodule41_not_fifomodule1), .Y(bouta_fifomodule41) );
	OR2X1 U2825 ( .A(bouta_fifomodule41), .B(boutb_fifomodule41), .Y(boutmain_fifomodule41) );
	DFFX2 U2826 ( .CLK(clk), .D(fifo_ocup_fifomodule41[0]), .Q(ocup_o[0]) );
	DFFX2 U2827 ( .CLK(clk), .D(fifo_ocup_fifomodule41[1]), .Q(ocup_o[1]) );
	DFFX2 U2828 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule41) );
	DFFX2 U2829 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule41) );
	DFFX2 U2830 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(write_ptr_ff_fifomodule41[0]) );
	DFFX2 U2831 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(read_ptr_ff_fifomodule41[0]) );
	DFFX2 U2832 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(fifo_ff_fifomodule41[0]) );
	DFFX2 U2833 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(write_ptr_ff_fifomodule41[1]) );
	DFFX2 U2834 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(read_ptr_ff_fifomodule41[1]) );
	DFFX2 U2835 ( .CLK(arst_value_fifomodule41), .D(1'b0), .Q(fifo_ff_fifomodule41[1]) );

	DFFX2 U2836 ( .CLK(clk), .D(next_write_ptr_fifomodule41[0]), .Q(write_ptr_ff_fifomodule41[0]) );
	DFFX2 U2837 ( .CLK(clk), .D(next_write_ptr_fifomodule41[1]), .Q(write_ptr_ff_fifomodule41[1]) );
	DFFX2 U2838 ( .CLK(clk), .D(next_read_ptr_fifomodule41[0]), .Q(read_ptr_ff_fifomodule41[0]) );
	DFFX2 U2839 ( .CLK(clk), .D(next_read_ptr_fifomodule41[1]), .Q(read_ptr_ff_fifomodule41[1]) );
	  

	DFFX2 U2840 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][0]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8]) );
	DFFX2 U2841 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][1]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+1]) );
	DFFX2 U2842 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][2]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+2]) );
	DFFX2 U2843 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][3]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+3]) );
	DFFX2 U2844 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][4]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+4]) );
	DFFX2 U2845 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][5]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+5]) );
	DFFX2 U2846 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][6]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+6]) );
	DFFX2 U2847 ( .CLK(u7temp_fifomodule41), .D(from_input_req_in_jump_input_datapath4put_datapath4[73:40][7]), .Q(fifo_ff_fifomodule41[write_ptr_ff_fifomodule41[0]*8+7]) );

    BUFX1 U2848 ( .A(locked_by_route_ff_vc_buffer41), .Y(next_locked_vc_buffer41) );
    BUFX1 U2849(.A(flit41[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][0]));
	BUFX1 U2850(.A(flit41[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][1]));
	BUFX1 U2851(.A(flit41[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][2]));
	BUFX1 U2852(.A(flit41[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][3]));
	BUFX1 U2853(.A(flit41[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][4]));
	BUFX1 U2854(.A(flit41[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][5]));
	BUFX1 U2855(.A(flit41[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][6]));
	BUFX1 U2856(.A(flit41[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][7]));
	BUFX1 U2857(.A(flit41[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][8]));
	BUFX1 U2858(.A(flit41[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][9]));
	BUFX1 U2859(.A(flit41[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][10]));
	BUFX1 U2860(.A(flit41[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][11]));
	BUFX1 U2861(.A(flit41[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][12]));
	BUFX1 U2862(.A(flit41[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][13]));
	BUFX1 U2863(.A(flit41[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][14]));
	BUFX1 U2864(.A(flit41[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][15]));
	BUFX1 U2865(.A(flit41[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][16]));
	BUFX1 U2866(.A(flit41[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][17]));
	BUFX1 U2867(.A(flit41[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][18]));
	BUFX1 U2868(.A(flit41[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][19]));
	BUFX1 U2869(.A(flit41[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][20]));
	BUFX1 U2870(.A(flit41[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][21]));
	BUFX1 U2871(.A(flit41[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][22]));
	BUFX1 U2872(.A(flit41[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][23]));
	BUFX1 U2873(.A(flit41[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][24]));
	BUFX1 U2874(.A(flit41[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][25]));
	BUFX1 U2875(.A(flit41[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][26]));
	BUFX1 U2876(.A(flit41[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][27]));
	BUFX1 U2877(.A(flit41[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][28]));
	BUFX1 U2878(.A(flit41[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][29]));
	BUFX1 U2879(.A(flit41[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][30]));
	BUFX1 U2880(.A(flit41[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][31]));
	BUFX1 U2881(.A(flit41[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][32]));
	BUFX1 U2882(.A(flit41[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[73:40][33]));
    NOR2X1 U2883 ( .IN1(flit41[33]), .IN2(flit41[32]), .QN(norres_vc_buffer41_vc_buffer1) );
    OR4X1 U2884 ( .IN1(flit41[29]), .IN2(flit41[28]), .IN3(flit41[27]), .IN4(flit41[26]), .Y(or1res_vc_buffer41) );
    OR4X1 U2885 ( .IN1(flit41[25]), .IN2(flit41[24]), .IN3(flit41[23]), .IN4(flit41[22]), .Y(or2res_vc_buffer41) );
    OR2X1 U2886 ( .A(or1res_vc_buffer41), .B(or2res_vc_buffer41), .Y(orres_vc_buffer41) );
    AND3X1 U2887 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(norres_vc_buffer41_vc_buffer1), .IN3(orres_vc_buffer41), .Q(finres1_vc_buffer41) );
    MUX21X1 U2888 (.IN1(next_locked_vc_buffer41), .IN2(1'b1), .S(finres1_vc_buffer41), .Q(next_locked_vc_buffer41);
    AND3X1 U2889 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(flit41[33]), .IN3(flit41[32]), .Q(andres1_vc_buffer41) );
    MUX21X1 U2890 (.IN1(next_locked_vc_buffer41), .IN2(1'b0), .S(andres1_vc_buffer41), .Q(next_locked_vc_buffer41);

    INVX1 U2891 ( .A(full_vc_buffer41), .Y(full_vc_buffer41_not1) );
    INVX1 U2892 ( .A(locked_by_route_ff_vc_buffer41), .Y(locked_by_route_ff_vc_buffer41_not1) );

    MUX21X1 U2893 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer41_not1), .S(norres_vc_buffer41_vc_buffer1), .Q(thirdand_vc_buffer41);
    AND3X1 U2894 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[37]), .IN2(full_vc_buffer41_not1), .IN3(thirdand_vc_buffer41), .Q(write_flit41_vc_buffer14) );
    AND2X1 U2895 ( .IN1(full_vc_buffer41_not1), .IN2(norres_vc_buffer41_vc_buffer1), .Q(from_input_resp_input_datapath4[1]) );
    INVX1 U2896 ( .A(empty_vc_buffer41), .Y(to_output_req_in_jump_input_datapath4put_datapath4[37]) );
    AND2X1 U2897 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[37]), .IN2(to_output_resp_input_datapath4[1]), .Q(read_flit41_vc_buffer14) );
	BUFX1 U2898(.A(to_output_req_in_jump_input_datapath4put_datapath4[39:38]), .Y(2'b01));

	DFFX2 U2899 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U2900 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U2901 (.IN1(next_locked_vc_buffer41), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer41);


	BUFX1 U2902 ( .A(read_ptr_ff_fifomodule42[0]), .Y(next_read_ptr_fifomodule42[0]) );
	BUFX1 U2903 ( .A(read_ptr_ff_fifomodule42[1]), .Y(next_read_ptr_fifomodule42[1]) );
	BUFX1 U2904 ( .A(write_ptr_ff_fifomodule42[0]), .Y(next_write_ptr_fifomodule42[0]) );
	BUFX1 U2905 ( .A(write_ptr_ff_fifomodule42[1]), .Y(next_write_ptr_fifomodule42[1]) );

	XNOR2X1 U2906 ( .IN1(write_ptr_ff_fifomodule42[0]), .IN2(read_ptr_ff_fifomodule42[0]), .Q(u1temp_fifomodule42) );
	XNOR2X1 U2907 ( .IN1(write_ptr_ff_fifomodule42[1]), .IN2(read_ptr_ff_fifomodule42[1]), .Q(u2temp_fifomodule42) );
	AND2X1 U2908 ( .A(u1temp_fifomodule42), .B(u2temp_fifomodule42), .Y(empty_vc_buffer42) );
	XOR2X1 U2909 ( .A(write_ptr_ff_fifomodule42[1]), .B(read_ptr_ff_fifomodule42[1]), .Y(u4temp_fifomodule42) );
	AND2X1 U2910 ( .A(u1temp_fifomodule42), .B(u4temp_fifomodule42), .Y(full_vc_buffer42) );
	MUX21X1 U2911 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][0]));
	MUX21X1 U2912 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+1]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][1]));
	MUX21X1 U2913 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+2]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][2]));
	MUX21X1 U2914 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+3]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][3]));
	MUX21X1 U2915 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+4]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][4]));
	MUX21X1 U2916 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+5]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][5]));
	MUX21X1 U2917 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+6]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][6]));
	MUX21X1 U2918 (.IN1(fifo_ff_fifomodule42[read_ptr_ff_fifomodule42[0] * 8+7]), .IN2(1'b0), .S(empty_vc_buffer42), .Q(to_output_req_in_jump_input_datapath4put_datapath4[110:77][7]));

	INVX1 U2919 ( .A(full_vc_buffer42), .Y(full_vc_buffer42_not2_fifomodule2) );
	AND2X1 U2920 ( .A(write_flit42_vc_buffer24), .B(full_vc_buffer42_not2_fifomodule2), .Y(u7temp_fifomodule42) );
	MUX21X1 U2921 (.IN1(1'b0), .IN2(1'b1), .S(u7temp_fifomodule42), .Q(u9temp_fifomodule42));
	HADDX1 U2922 ( .A0(write_ptr_ff_fifomodule42[0]), .B0(u9temp_fifomodule42), .C1(u10carry_fifomodule42), .SO(next_write_ptr_fifomodule42[0]) );
	HADDX1 U2923 ( .A0(u10carry_fifomodule42), .B0(write_ptr_ff_fifomodule42[1]), .C1(u11carry_fifomodule42), .SO(next_write_ptr_fifomodule42[1]) );

	INVX1 U2924 ( .A(empty_vc_buffer42), .Y(empty_vc_buffer42_not_fifomodule2) );
	AND2X1 U2925 ( .A(read_flit42_vc_buffer24), .B(empty_vc_buffer42_not_fifomodule2), .Y(u13temp_fifomodule42) );
	MUX21X1 U2926 (.IN1(1'b0), .IN2(1'b1), .S(u13temp_fifomodule42), .Q(u14temp_fifomodule42));
	HADDX1 U2927 ( .A0(read_ptr_ff_fifomodule42[0]), .B0(u14temp_fifomodule42), .C1(u15carry_fifomodule42), .SO(next_read_ptr_fifomodule42[0]) );
	HADDX1 U2928 ( .A0(u15carry_fifomodule42), .B0(read_ptr_ff_fifomodule42[1]), .C1(u16carry_fifomodule42), .SO(next_read_ptr_fifomodule42[1]) );

	AND2X1 U2929 ( .A(write_flit42_vc_buffer24), .B(full_vc_buffer42), .Y(u17res_fifomodule42) );
	AND2X1 U2930 ( .A(read_flit42_vc_buffer24), .B(empty_vc_buffer42), .Y(u18res_fifomodule42) );
    OR2X1 U2931 ( .A(u17res_fifomodule42), .B(u18res_fifomodule42), .Y(error_vc_buffer42) );
	XOR2X1 U2932 ( .A(write_ptr_ff_fifomodule42[0]), .B(read_ptr_ff_fifomodule42[0]), .Y(fifo_ocup_fifomodule42[0]) );
	INVX1 U2933 ( .A(write_ptr_ff_fifomodule42[0]), .Y(write_ptr_ff_fifomodule42_0_not24) );
	AND2X1 U2934 ( .A(write_ptr_ff_fifomodule42_0_not24), .B(read_ptr_ff_fifomodule42[0]), .Y(b0wire_fifomodule42) );
	XOR2X1 U2935 ( .A(write_ptr_ff_fifomodule42[1]), .B(read_ptr_ff_fifomodule42[1]), .Y(u23temp_fifomodule42) );
	INVX1 U2936 ( .A(write_ptr_ff_fifomodule42[1]), .Y(write_ptr_ff_fifomodule42_1_not24) );
	AND2X1 U2937 ( .A(read_ptr_ff_fifomodule42[1]), .B(write_ptr_ff_fifomodule42_1_not24), .Y(boutb_fifomodule42) );
	XOR2X1 U2938 ( .A(u23temp_fifomodule42), .B(b0wire_fifomodule42), .Y(fifo_ocup_fifomodule42[1]) );
	INVX1 U2939 ( .A(u23temp_fifomodule42), .Y(u23temp_fifomodule42_not_fifomodule2) );
	AND2X1 U2940 ( .A(b0wire_fifomodule42), .B(u23temp_fifomodule42_not_fifomodule2), .Y(bouta_fifomodule42) );
	OR2X1 U2941 ( .A(bouta_fifomodule42), .B(boutb_fifomodule42), .Y(boutmain_fifomodule42) );
	DFFX2 U2942 ( .CLK(clk), .D(fifo_ocup_fifomodule42[0]), .Q(ocup_o[0]) );
	DFFX2 U2943 ( .CLK(clk), .D(fifo_ocup_fifomodule42[1]), .Q(ocup_o[1]) );
	DFFX2 U2944 ( .CLK(clk), .D(arst), .Q(arst_value_fifomodule42) );
	DFFX2 U2945 ( .CLK(arst), .D(arst), .Q(arst_value_fifomodule42) );
	DFFX2 U2946 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(write_ptr_ff_fifomodule42[0]) );
	DFFX2 U2947 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(read_ptr_ff_fifomodule42[0]) );
	DFFX2 U2948 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(fifo_ff_fifomodule42[0]) );
	DFFX2 U2949 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(write_ptr_ff_fifomodule42[1]) );
	DFFX2 U2950 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(read_ptr_ff_fifomodule42[1]) );
	DFFX2 U2951 ( .CLK(arst_value_fifomodule42), .D(1'b0), .Q(fifo_ff_fifomodule42[1]) );

	DFFX2 U2952 ( .CLK(clk), .D(next_write_ptr_fifomodule42[0]), .Q(write_ptr_ff_fifomodule42[0]) );
	DFFX2 U2953 ( .CLK(clk), .D(next_write_ptr_fifomodule42[1]), .Q(write_ptr_ff_fifomodule42[1]) );
	DFFX2 U2954 ( .CLK(clk), .D(next_read_ptr_fifomodule42[0]), .Q(read_ptr_ff_fifomodule42[0]) );
	DFFX2 U2955 ( .CLK(clk), .D(next_read_ptr_fifomodule42[1]), .Q(read_ptr_ff_fifomodule42[1]) );
	  

	DFFX2 U2956 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][0]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8]) );
	DFFX2 U2957 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][1]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+1]) );
	DFFX2 U2958 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][2]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+2]) );
	DFFX2 U2959 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][3]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+3]) );
	DFFX2 U2960 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][4]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+4]) );
	DFFX2 U2961 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][5]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+5]) );
	DFFX2 U2962 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][6]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+6]) );
	DFFX2 U2963 ( .CLK(u7temp_fifomodule42), .D(from_input_req_in_jump_input_datapath4put_datapath4[110:77][7]), .Q(fifo_ff_fifomodule42[write_ptr_ff_fifomodule42[0]*8+7]) );

    BUFX1 U2964 ( .A(locked_by_route_ff_vc_buffer42), .Y(next_locked_vc_buffer42) );
    BUFX1 U2965(.A(flit42[0]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][0]));
	BUFX1 U2966(.A(flit42[1]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][1]));
	BUFX1 U2967(.A(flit42[2]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][2]));
	BUFX1 U2968(.A(flit42[3]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][3]));
	BUFX1 U2969(.A(flit42[4]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][4]));
	BUFX1 U2970(.A(flit42[5]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][5]));
	BUFX1 U2971(.A(flit42[6]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][6]));
	BUFX1 U2972(.A(flit42[7]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][7]));
	BUFX1 U2973(.A(flit42[8]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][8]));
	BUFX1 U2974(.A(flit42[9]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][9]));
	BUFX1 U2975(.A(flit42[10]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][10]));
	BUFX1 U2976(.A(flit42[11]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][11]));
	BUFX1 U2977(.A(flit42[12]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][12]));
	BUFX1 U2978(.A(flit42[13]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][13]));
	BUFX1 U2979(.A(flit42[14]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][14]));
	BUFX1 U2980(.A(flit42[15]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][15]));
	BUFX1 U2981(.A(flit42[16]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][16]));
	BUFX1 U2982(.A(flit42[17]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][17]));
	BUFX1 U2983(.A(flit42[18]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][18]));
	BUFX1 U2984(.A(flit42[19]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][19]));
	BUFX1 U2985(.A(flit42[20]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][20]));
	BUFX1 U2986(.A(flit42[21]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][21]));
	BUFX1 U2987(.A(flit42[22]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][22]));
	BUFX1 U2988(.A(flit42[23]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][23]));
	BUFX1 U2989(.A(flit42[24]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][24]));
	BUFX1 U2990(.A(flit42[25]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][25]));
	BUFX1 U2991(.A(flit42[26]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][26]));
	BUFX1 U2992(.A(flit42[27]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][27]));
	BUFX1 U2993(.A(flit42[28]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][28]));
	BUFX1 U2994(.A(flit42[29]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][29]));
	BUFX1 U2995(.A(flit42[30]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][30]));
	BUFX1 U2996(.A(flit42[31]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][31]));
	BUFX1 U2997(.A(flit42[32]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][32]));
	BUFX1 U2998(.A(flit42[33]), .Y(from_input_req_in_jump_input_datapath4put_datapath4[110:77][33]));
    NOR2X1 U2999 ( .IN1(flit42[33]), .IN2(flit42[32]), .QN(norres_vc_buffer42_vc_buffer2) );
    OR4X1 U3000 ( .IN1(flit42[29]), .IN2(flit42[28]), .IN3(flit42[27]), .IN4(flit42[26]), .Y(or1res_vc_buffer42) );
    OR4X1 U3001 ( .IN1(flit42[25]), .IN2(flit42[24]), .IN3(flit42[23]), .IN4(flit42[22]), .Y(or2res_vc_buffer42) );
    OR2X1 U3002 ( .A(or1res_vc_buffer42), .B(or2res_vc_buffer42), .Y(orres_vc_buffer42) );
    AND3X1 U3003 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(norres_vc_buffer42_vc_buffer2), .IN3(orres_vc_buffer42), .Q(finres1_vc_buffer42) );
    MUX21X1 U3004 (.IN1(next_locked_vc_buffer42), .IN2(1'b1), .S(finres1_vc_buffer42), .Q(next_locked_vc_buffer42);
    AND3X1 U3005 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(flit42[33]), .IN3(flit42[32]), .Q(andres1_vc_buffer42) );
    MUX21X1 U3006 (.IN1(next_locked_vc_buffer42), .IN2(1'b0), .S(andres1_vc_buffer42), .Q(next_locked_vc_buffer42);

    INVX1 U3007 ( .A(full_vc_buffer42), .Y(full_vc_buffer42_not2) );
    INVX1 U3008 ( .A(locked_by_route_ff_vc_buffer42), .Y(locked_by_route_ff_vc_buffer42_not2) );

    MUX21X1 U3009 (.IN1(1'b1), .IN2(locked_by_route_ff_vc_buffer42_not2), .S(norres_vc_buffer42_vc_buffer2), .Q(thirdand_vc_buffer42);
    AND3X1 U3010 ( .IN1(from_input_req_in_jump_input_datapath4put_datapath4[74]), .IN2(full_vc_buffer42_not2), .IN3(thirdand_vc_buffer42), .Q(write_flit42_vc_buffer24) );
    AND2X1 U3011 ( .IN1(full_vc_buffer42_not2), .IN2(norres_vc_buffer42_vc_buffer2), .Q(from_input_resp_input_datapath4[2]) );
    INVX1 U3012 ( .A(empty_vc_buffer42), .Y(to_output_req_in_jump_input_datapath4put_datapath4[74]) );
    AND2X1 U3013 ( .IN1(to_output_req_in_jump_input_datapath4put_datapath4[74]), .IN2(to_output_resp_input_datapath4[2]), .Q(read_flit42_vc_buffer24) );
	BUFX1 U3014(.A(to_output_req_in_jump_input_datapath4put_datapath4[76:75]), .Y(2'b10));

	DFFX2 U3015 ( .CLK(clk), .D(arst), .Q(arst_value) );
    DFFX2 U3016 ( .CLK(arst), .D(arst), .Q(arst_value) );
    MUX21X1 U3017 (.IN1(next_locked_vc_buffer42), .IN2(1'sb0), .S(arst_value), .Q(locked_by_route_ff_vc_buffer42);

	BUFX1 U3018(.A(from_input_req_in_jump_input_datapath4put_datapath4[77]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U3019(.A(from_input_req_in_jump_input_datapath4put_datapath4[78]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U3020(.A(from_input_req_in_jump_input_datapath4put_datapath4[79]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U3021(.A(from_input_req_in_jump_input_datapath4put_datapath4[80]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U3022(.A(from_input_req_in_jump_input_datapath4put_datapath4[81]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U3023(.A(from_input_req_in_jump_input_datapath4put_datapath4[82]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U3024(.A(from_input_req_in_jump_input_datapath4put_datapath4[83]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U3025(.A(from_input_req_in_jump_input_datapath4put_datapath4[84]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U3026(.A(from_input_req_in_jump_input_datapath4put_datapath4[85]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U3027(.A(from_input_req_in_jump_input_datapath4put_datapath4[86]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U3028(.A(from_input_req_in_jump_input_datapath4put_datapath4[87]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U3029(.A(from_input_req_in_jump_input_datapath4put_datapath4[88]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U3030(.A(from_input_req_in_jump_input_datapath4put_datapath4[89]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U3031(.A(from_input_req_in_jump_input_datapath4put_datapath4[90]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U3032(.A(from_input_req_in_jump_input_datapath4put_datapath4[91]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U3033(.A(from_input_req_in_jump_input_datapath4put_datapath4[92]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U3034(.A(from_input_req_in_jump_input_datapath4put_datapath4[93]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U3035(.A(from_input_req_in_jump_input_datapath4put_datapath4[94]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U3036(.A(from_input_req_in_jump_input_datapath4put_datapath4[95]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U3037(.A(from_input_req_in_jump_input_datapath4put_datapath4[96]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U3038(.A(from_input_req_in_jump_input_datapath4put_datapath4[97]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U3039(.A(from_input_req_in_jump_input_datapath4put_datapath4[98]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U3040(.A(from_input_req_in_jump_input_datapath4put_datapath4[99]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U3041(.A(from_input_req_in_jump_input_datapath4put_datapath4[100]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U3042(.A(from_input_req_in_jump_input_datapath4put_datapath4[101]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U3043(.A(from_input_req_in_jump_input_datapath4put_datapath4[102]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U3044(.A(from_input_req_in_jump_input_datapath4put_datapath4[103]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U3045(.A(from_input_req_in_jump_input_datapath4put_datapath4[104]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U3046(.A(from_input_req_in_jump_input_datapath4put_datapath4[105]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U3047(.A(from_input_req_in_jump_input_datapath4put_datapath4[106]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U3048(.A(from_input_req_in_jump_input_datapath4put_datapath4[107]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U3049(.A(from_input_req_in_jump_input_datapath4put_datapath4[108]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U3050(.A(from_input_req_in_jump_input_datapath4put_datapath4[109]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U3051(.A(from_input_req_in_jump_input_datapath4put_datapath4[110]), .Y(ext_req_v_i[184:148][36]));
    XNOR2X1 U3052 ( .IN1(ext_req_v_i[184:148][1]), .IN2(i_input_datapath4[0]), .QN(xnor1resu_input_datapath4) );
    XNOR2X1 U3053 ( .IN1(ext_req_v_i[184:148][2]), .IN2(i_input_datapath4[1]), .QN(xnor2resu_input_datapath4) );
    AND2X1 U3054 ( .IN1(xnor1resu_input_datapath4), .IN2(xnor2resu_input_datapath4), .Q(and1resu_input_datapath4) );
    AND3X1 U3055 ( .IN1(and1resu_input_datapath4), .IN2(ext_req_v_i[184:148][0]), .IN2(ext_req_v_i[184:148][0]), .Q(cond1line_input_datapath4) );
    MUX21X1 U3056 (.IN1(vc_ch_act_in_input_datapath4[0]), .IN2(i_input_datapath4[0]), .S(cond1line_input_datapath4), .Q(vc_ch_act_in_input_datapath4[0]));
    MUX21X1 U3057 (.IN1(vc_ch_act_in_input_datapath4[1]), .IN2(i_input_datapath4[1]), .S(cond1line_input_datapath4), .Q(vc_ch_act_in_input_datapath4[1]));
    MUX21X1 U3058 (.IN1(req_in_jump_input_datapath4), .IN2(1), .S(cond1line_input_datapath4), .Q(req_in_jump_input_datapath4));
	BUFX1 U3059(.A(from_input_req_in_jump_input_datapath4put_datapath4[40]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U3060(.A(from_input_req_in_jump_input_datapath4put_datapath4[41]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U3061(.A(from_input_req_in_jump_input_datapath4put_datapath4[42]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U3062(.A(from_input_req_in_jump_input_datapath4put_datapath4[43]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U3063(.A(from_input_req_in_jump_input_datapath4put_datapath4[44]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U3064(.A(from_input_req_in_jump_input_datapath4put_datapath4[45]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U3065(.A(from_input_req_in_jump_input_datapath4put_datapath4[46]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U3066(.A(from_input_req_in_jump_input_datapath4put_datapath4[47]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U3067(.A(from_input_req_in_jump_input_datapath4put_datapath4[48]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U3068(.A(from_input_req_in_jump_input_datapath4put_datapath4[49]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U3069(.A(from_input_req_in_jump_input_datapath4put_datapath4[50]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U3070(.A(from_input_req_in_jump_input_datapath4put_datapath4[51]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U3071(.A(from_input_req_in_jump_input_datapath4put_datapath4[52]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U3072(.A(from_input_req_in_jump_input_datapath4put_datapath4[53]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U3073(.A(from_input_req_in_jump_input_datapath4put_datapath4[54]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U3074(.A(from_input_req_in_jump_input_datapath4put_datapath4[55]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U3075(.A(from_input_req_in_jump_input_datapath4put_datapath4[56]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U3076(.A(from_input_req_in_jump_input_datapath4put_datapath4[57]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U3077(.A(from_input_req_in_jump_input_datapath4put_datapath4[58]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U3078(.A(from_input_req_in_jump_input_datapath4put_datapath4[59]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U3079(.A(from_input_req_in_jump_input_datapath4put_datapath4[60]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U3080(.A(from_input_req_in_jump_input_datapath4put_datapath4[61]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U3081(.A(from_input_req_in_jump_input_datapath4put_datapath4[62]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U3082(.A(from_input_req_in_jump_input_datapath4put_datapath4[63]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U3083(.A(from_input_req_in_jump_input_datapath4put_datapath4[64]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U3084(.A(from_input_req_in_jump_input_datapath4put_datapath4[65]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U3085(.A(from_input_req_in_jump_input_datapath4put_datapath4[66]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U3086(.A(from_input_req_in_jump_input_datapath4put_datapath4[67]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U3087(.A(from_input_req_in_jump_input_datapath4put_datapath4[68]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U3088(.A(from_input_req_in_jump_input_datapath4put_datapath4[69]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U3089(.A(from_input_req_in_jump_input_datapath4put_datapath4[70]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U3090(.A(from_input_req_in_jump_input_datapath4put_datapath4[71]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U3091(.A(from_input_req_in_jump_input_datapath4put_datapath4[72]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U3092(.A(from_input_req_in_jump_input_datapath4put_datapath4[73]), .Y(ext_req_v_i[184:148][36]));

	BUFX1 U3093(.A(from_input_req_in_jump_input_datapath4put_datapath4[3]), .Y(ext_req_v_i[184:148][3]));
	BUFX1 U3094(.A(from_input_req_in_jump_input_datapath4put_datapath4[4]), .Y(ext_req_v_i[184:148][4]));
	BUFX1 U3095(.A(from_input_req_in_jump_input_datapath4put_datapath4[5]), .Y(ext_req_v_i[184:148][5]));
	BUFX1 U3096(.A(from_input_req_in_jump_input_datapath4put_datapath4[6]), .Y(ext_req_v_i[184:148][6]));
	BUFX1 U3097(.A(from_input_req_in_jump_input_datapath4put_datapath4[7]), .Y(ext_req_v_i[184:148][7]));
	BUFX1 U3098(.A(from_input_req_in_jump_input_datapath4put_datapath4[8]), .Y(ext_req_v_i[184:148][8]));
	BUFX1 U3099(.A(from_input_req_in_jump_input_datapath4put_datapath4[9]), .Y(ext_req_v_i[184:148][9]));
	BUFX1 U3100(.A(from_input_req_in_jump_input_datapath4put_datapath4[10]), .Y(ext_req_v_i[184:148][10]));
	BUFX1 U3101(.A(from_input_req_in_jump_input_datapath4put_datapath4[11]), .Y(ext_req_v_i[184:148][11]));
	BUFX1 U3102(.A(from_input_req_in_jump_input_datapath4put_datapath4[12]), .Y(ext_req_v_i[184:148][12]));
	BUFX1 U3103(.A(from_input_req_in_jump_input_datapath4put_datapath4[13]), .Y(ext_req_v_i[184:148][13]));
	BUFX1 U3104(.A(from_input_req_in_jump_input_datapath4put_datapath4[14]), .Y(ext_req_v_i[184:148][14]));
	BUFX1 U3105(.A(from_input_req_in_jump_input_datapath4put_datapath4[15]), .Y(ext_req_v_i[184:148][15]));
	BUFX1 U3106(.A(from_input_req_in_jump_input_datapath4put_datapath4[16]), .Y(ext_req_v_i[184:148][16]));
	BUFX1 U3107(.A(from_input_req_in_jump_input_datapath4put_datapath4[17]), .Y(ext_req_v_i[184:148][17]));
	BUFX1 U3108(.A(from_input_req_in_jump_input_datapath4put_datapath4[18]), .Y(ext_req_v_i[184:148][18]));
	BUFX1 U3109(.A(from_input_req_in_jump_input_datapath4put_datapath4[19]), .Y(ext_req_v_i[184:148][19]));
	BUFX1 U3110(.A(from_input_req_in_jump_input_datapath4put_datapath4[20]), .Y(ext_req_v_i[184:148][20]));
	BUFX1 U3111(.A(from_input_req_in_jump_input_datapath4put_datapath4[21]), .Y(ext_req_v_i[184:148][21]));
	BUFX1 U3112(.A(from_input_req_in_jump_input_datapath4put_datapath4[22]), .Y(ext_req_v_i[184:148][22]));
	BUFX1 U3113(.A(from_input_req_in_jump_input_datapath4put_datapath4[23]), .Y(ext_req_v_i[184:148][23]));
	BUFX1 U3114(.A(from_input_req_in_jump_input_datapath4put_datapath4[24]), .Y(ext_req_v_i[184:148][24]));
	BUFX1 U3115(.A(from_input_req_in_jump_input_datapath4put_datapath4[25]), .Y(ext_req_v_i[184:148][25]));
	BUFX1 U3116(.A(from_input_req_in_jump_input_datapath4put_datapath4[26]), .Y(ext_req_v_i[184:148][26]));
	BUFX1 U3117(.A(from_input_req_in_jump_input_datapath4put_datapath4[27]), .Y(ext_req_v_i[184:148][27]));
	BUFX1 U3118(.A(from_input_req_in_jump_input_datapath4put_datapath4[28]), .Y(ext_req_v_i[184:148][28]));
	BUFX1 U3119(.A(from_input_req_in_jump_input_datapath4put_datapath4[29]), .Y(ext_req_v_i[184:148][29]));
	BUFX1 U3120(.A(from_input_req_in_jump_input_datapath4put_datapath4[30]), .Y(ext_req_v_i[184:148][30]));
	BUFX1 U3121(.A(from_input_req_in_jump_input_datapath4put_datapath4[31]), .Y(ext_req_v_i[184:148][31]));
	BUFX1 U3122(.A(from_input_req_in_jump_input_datapath4put_datapath4[32]), .Y(ext_req_v_i[184:148][32]));
	BUFX1 U3123(.A(from_input_req_in_jump_input_datapath4put_datapath4[33]), .Y(ext_req_v_i[184:148][33]));
	BUFX1 U3124(.A(from_input_req_in_jump_input_datapath4put_datapath4[34]), .Y(ext_req_v_i[184:148][34]));
	BUFX1 U3125(.A(from_input_req_in_jump_input_datapath4put_datapath4[35]), .Y(ext_req_v_i[184:148][35]));
	BUFX1 U3126(.A(from_input_req_in_jump_input_datapath4put_datapath4[36]), .Y(ext_req_v_i[184:148][36]));

    MUX21X1 U3127 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4 * 37]), .IN2(ext_req_v_i[184:148][0]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4 * 37]));
    MUX21X1 U3128 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+2]), .IN2(vc_ch_act_in_input_datapath4[1]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+2]));
    MUX21X1 U3129 (.IN1(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+1]), .IN2(vc_ch_act_in_input_datapath4[0]), .S(req_in_jump_input_datapath4), .Q(from_input_req_in_jump_input_datapath4put_datapath4[vc_ch_act_in_input_datapath4*37+1]));
    MUX21X1 U3130 (.IN1(ext_resp_v_o[5:4][0]), .IN2(from_input_resp_input_datapath4[vc_ch_act_in_input_datapath4]), .S(req_in_jump_input_datapath4), .Q(ext_resp_v_o[5:4][0]));

    INVX1 U3131 ( .A(req_in_jump_input_datapath4), .Y(req_in_jump_input_datapath4_not) );
    MUX21X1 U3132 (.IN1(ext_resp_v_o[5:4][0]), .IN2(1'sb1), .S(req_in_jump_input_datapath4_not), .Q(ext_resp_v_o[5:4][0]));
    BUFX1 U3133(.A(from_input_req_in_jump_input_datapath4put_datapath4[34]), .Y(ext_req_v_i[184:148][34]));

    XOR2X1 U3134 ( .IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b1), .Q(xor1resu_input_datapath4) );
    MUX21X1 U3135 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(xor1resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U3136 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b0), .S(xor1resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[1]));
    AND2X1 U3137 ( .IN1(xor1resu_input_datapath4), .IN2(to_output_req_in_jump_input_datapath4put_datapath4[j_input_datapath4*37]), .Q(and2resu_input_datapath4) );
    MUX21X1 U3138 (.IN1(vc_ch_act_out_input_datapath4[0]), .IN2(j_input_datapath4[0]), .S(and2resu_input_datapath4), .Q(vc_ch_act_out_input_datapath4[0]));
    MUX21X1 U3139 (.IN1(vc_ch_act_out_input_datapath4[1]), .IN2(j_input_datapath4[1]), .S(and2resu_input_datapath4), .Q(vc_ch_act_out_input_datapath4[1]));
    MUX21X1 U3140 (.IN1(req_out_jump_input_datapath4), .IN2(1'b1), .S(and2resu_input_datapath4), .Q(req_out_jump_input_datapath4));
    MUX21X1 U3141 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(and2resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U3142 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b1), .S(and2resu_input_datapath4), .Q(_sv2v_jump_input_datapath4[1]));
    HADDX1 U3143 ( .A0(j_input_datapath4[0]), .B0(1'b1), .C1(j_input_datapath4[1]), .SO(j_input_datapath4[0]) );
    HADDX1 U3144 ( .A0(j_input_datapath4[0]), .B0(1'b1), .C1(j_input_datapath4[1]), .SO(j_input_datapath4[0]) );
    AND2X1 U3145 ( .IN1(xor1resu_input_datapath4), .IN2(to_output_req_in_jump_input_datapath4put_datapath4[j_input_datapath4*37]), .Q(and3resu) );
    NAND2X1 U3146(.A(_sv2v_jump_input_datapath4[0]),.B(_sv2v_jump_input_datapath4[1]),.Y(nand1resu_input_datapath44));
    MUX21X1 U3147 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(1'b0), .S(nand1resu_input_datapath44), .Q(_sv2v_jump_input_datapath4[0]));
    MUX21X1 U3148 (.IN1(_sv2v_jump_input_datapath4[1]), .IN2(1'b0), .S(nand1resu_input_datapath44), .Q(_sv2v_jump_input_datapath4[1]));
    XNOR2X1 U3149 (.IN1(_sv2v_jump_input_datapath4[0]), .IN2(_sv2v_jump_input_datapath4[1]), .Q(xnor23resu_input_datapath4) );
    AND2X1 U3150 ( .IN1(xnor23resu_input_datapath4), .IN2(req_out_jump_input_datapath4), .Q(and4resu_input_datapath4) );

    MUX21X1 U3151(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+3]),.IN2(int_req_v[184:148][3]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+3]));
	MUX21X1 U3152(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+4]),.IN2(int_req_v[184:148][4]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+4]));
	MUX21X1 U3153(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+5]),.IN2(int_req_v[184:148][5]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+5]));
	MUX21X1 U3154(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+6]),.IN2(int_req_v[184:148][6]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+6]));
	MUX21X1 U3155(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+7]),.IN2(int_req_v[184:148][7]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+7]));
	MUX21X1 U3156(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+8]),.IN2(int_req_v[184:148][8]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+8]));
	MUX21X1 U3157(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+9]),.IN2(int_req_v[184:148][9]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+9]));
	MUX21X1 U3158(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+10]),.IN2(int_req_v[184:148][10]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+10]));
	MUX21X1 U3159(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+11]),.IN2(int_req_v[184:148][11]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+11]));
	MUX21X1 U3160(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+12]),.IN2(int_req_v[184:148][12]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+12]));
	MUX21X1 U3161(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+13]),.IN2(int_req_v[184:148][13]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+13]));
	MUX21X1 U3162(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+14]),.IN2(int_req_v[184:148][14]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+14]));
	MUX21X1 U3163(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+15]),.IN2(int_req_v[184:148][15]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+15]));
	MUX21X1 U3164(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+16]),.IN2(int_req_v[184:148][16]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+16]));
	MUX21X1 U3165(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+17]),.IN2(int_req_v[184:148][17]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+17]));
	MUX21X1 U3166(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+18]),.IN2(int_req_v[184:148][18]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+18]));
	MUX21X1 U3167(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+19]),.IN2(int_req_v[184:148][19]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+19]));
	MUX21X1 U3168(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+20]),.IN2(int_req_v[184:148][20]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+20]));
	MUX21X1 U3169(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+21]),.IN2(int_req_v[184:148][21]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+21]));
	MUX21X1 U3170(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+22]),.IN2(int_req_v[184:148][22]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+22]));
	MUX21X1 U3171(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+23]),.IN2(int_req_v[184:148][23]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+23]));
	MUX21X1 U3172(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+24]),.IN2(int_req_v[184:148][24]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+24]));
	MUX21X1 U3173(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+25]),.IN2(int_req_v[184:148][25]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+25]));
	MUX21X1 U3174(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+26]),.IN2(int_req_v[184:148][26]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+26]));
	MUX21X1 U3175(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+27]),.IN2(int_req_v[184:148][27]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+27]));
	MUX21X1 U3176(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+28]),.IN2(int_req_v[184:148][28]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+28]));
	MUX21X1 U3177(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+29]),.IN2(int_req_v[184:148][29]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+29]));
	MUX21X1 U3178(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+30]),.IN2(int_req_v[184:148][30]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+30]));
	MUX21X1 U3179(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+31]),.IN2(int_req_v[184:148][31]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+31]));
	MUX21X1 U3180(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+32]),.IN2(int_req_v[184:148][32]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+32]));
	MUX21X1 U3181(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+33]),.IN2(int_req_v[184:148][33]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+33]));
	MUX21X1 U3182(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+34]),.IN2(int_req_v[184:148][34]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+34]));
	MUX21X1 U3183(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+35]),.IN2(int_req_v[184:148][35]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+35]));
	MUX21X1 U3184(.IN1(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+36]),.IN2(int_req_v[184:148][36]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_ouot*37)+36]));

	MUX21X1 U3185(.IN1(int_req_v[184:148][0]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4 * 37)]), .S(and4resu_input_datapath4), .Q(int_req_v[184:148][0]));
	MUX21X1 U3186(.IN1(int_req_v[184:148][1]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+1]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+1]));
	MUX21X1 U3187(.IN1(int_req_v[184:148][2]),.IN2(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+2]), .S(and4resu_input_datapath4), .Q(to_output_req_in_jump_input_datapath4put_datapath4[(vc_ch_act_out_input_datapath4*37)+2]));
	MUX21X1 U3188(.IN1(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4]),.IN2(int_resp_v[5:4]), .S(and4resu_input_datapath4), .Q(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4]));
	MUX21X1 U3189(.IN1(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4+1]),.IN2(int_resp_v[5:4]), .S(and4resu_input_datapath4), .Q(to_output_resp_input_datapath4[vc_ch_act_out_input_datapath4+1]));



//output part	

    BUFX1 U3190 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[0]) );
    BUFX1 U3191 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1[1]) );
    BUFX1 U3192 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3193 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3194 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    XNOR2X1 U3195 ( .IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1) );
    MUX21X1 U3196 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U3197 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    INVX1 U3198 ( .A(i_high_prior_arbiter1[0]), .Y(i_0_not_high_prior_arbiter1) );
    MUX21X1 U3199 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[0]);
    MUX21X1 U3200 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1[0]), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(raw_grant[1]);
    MUX21X1 U3201 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U3202 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b1), .S(valid_from_im_output_module[3:0][i_high_prior_arbiter1[0]]), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    NAND2X1 U3203 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(_sv2v_jump_high_prior_arbiter1[1]), .QN(nandres_high_prior_arbiter1) );
    MUX21X1 U3204 (.IN1(_sv2v_jump_high_prior_arbiter1[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[0]));
    MUX21X1 U3205 (.IN1(_sv2v_jump_high_prior_arbiter1[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1), .Q(_sv2v_jump_high_prior_arbiter1[1]));
    HADDX1 U3206 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U3207 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );
    HADDX1 U3208 ( .A0(i_high_prior_arbiter1[0]), .B0(1'b1), .C1(i_high_prior_arbiter1[1]), .SO(i_high_prior_arbiter1[0]) );



    BUFX1 U3209 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[0]) );
    BUFX1 U3210 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2[1]) );
    BUFX1 U3211 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3212 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3213 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    XNOR2X1 U3214 ( .IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2) );
    MUX21X1 U3215 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U3216 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    INVX1 U3217 ( .A(i_high_prior_arbiter2[0]), .Y(i_0_not_high_prior_arbiter2) );
    MUX21X1 U3218 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[0]);
    MUX21X1 U3219 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2[0]), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(masked_grant[1]);
    MUX21X1 U3220 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U3221 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2[0]]), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    NAND2X1 U3222 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(_sv2v_jump_high_prior_arbiter2[1]), .QN(nandres_high_prior_arbiter2) );
    MUX21X1 U3223 (.IN1(_sv2v_jump_high_prior_arbiter2[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[0]));
    MUX21X1 U3224 (.IN1(_sv2v_jump_high_prior_arbiter2[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2), .Q(_sv2v_jump_high_prior_arbiter2[1]));
    HADDX1 U3225 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U3226 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    HADDX1 U3227 ( .A0(i_high_prior_arbiter2[0]), .B0(1'b1), .C1(i_high_prior_arbiter2[1]), .SO(i_high_prior_arbiter2[0]) );
    

    BUFX1 U3228 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[0]) );
    BUFX1 U3229 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter[1]) );
    AND2X1 U3230 ( .A(mask_ff_rr_arbiter[0]), .B(valid_from_im_output_module[3:0][0]), .Y(mask_req_rr_arbiter[0]) );
    AND2X1 U3231 ( .A(mask_ff_rr_arbiter[1]), .B(valid_from_im_output_module[3:0][1]), .Y(mask_req_rr_arbiter[1]) );
    BUFX1 U3232 ( .A(mask_ff_rr_arbiter[0]), .Y(next_mask_rr_arbiter[0]) );
    BUFX1 U3233 ( .A(mask_ff_rr_arbiter[1]), .Y(next_mask_rr_arbiter[1]) );
    XNOR2X1 U3234 ( .IN1(mask_req_rr_arbiter[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter) );
    XNOR2X1 U3235 ( .IN1(mask_req_rr_arbiter[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter) );
    MUX21X1 U3236 (.IN1(masked_grant_rr_arbiter[0]), .IN2(raw_grant_rr_arbiter[0]), .S(xnor0res_rr_arbiter), .Q(grant_im_output_module[3:0][0]));
    MUX21X1 U3237 (.IN1(masked_grant_rr_arbiter[1]), .IN2(raw_grant_rr_arbiter[1]), .S(xnor1res_rr_arbiter), .Q(grant_im_output_module[3:0][1]));

    BUFX1 U3238 ( .A(1'b0), .Y(i_rr_arbiter[1]) );
    MUX21X1 U3239 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter[0]));

    AND2X1 U3240 ( .A(_sv2v_jump_rr_rr_arbiter[1]), .B(1'b0), .Y(firstif_rr_arbiter) );
    MUX21X1 U3241 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U3242 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(firstif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    AND2X1 U3243 ( .A(firstif_rr_arbiter), .B(grant_im_output_module[3:0][i_rr_arbiter[0]]), .Y(secondif_rr_arbiter) );
    MUX21X1 U3244 (.IN1(next_mask_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[0]));
    MUX21X1 U3245 (.IN1(next_mask_rr_arbiter[1]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(next_mask_rr_arbiter[1]));
    MUX21X1 U3246 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter[0]), .Q(j_rr_arbiter[0]));
    AND2X1 U3247 ( .A(secondif_rr_arbiter), .B(j_rr_arbiter[0]), .Y(thirdif_rr_arbiter) );
    MUX21X1 U3248 (.IN1(next_mask_rr_arbiter[j_rr_arbiter[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter), .Q(next_mask_rr_arbiter[j_rr_arbiter[0]]));
    MUX21X1 U3249 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U3250 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b1), .S(secondif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));
    NAND2X1 U3251 ( .IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(_sv2v_jump_rr_rr_arbiter[1]), .QN(fourthif_rr_arbiter) );
    MUX21X1 U3252 (.IN1(_sv2v_jump_rr_rr_arbiter[0]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[0]));
    MUX21X1 U3253 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(fourthif_rr_arbiter), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    MUX21X1 U3254 (.IN1(_sv2v_jump_rr_rr_arbiter[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter[1]));

    DFFX2 U3255 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter) );
    DFFX2 U3256 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter) );
    MUX21X1 U3257 (.IN1(mask_ff_rr_arbiter[0]), .IN2(next_mask_rr_arbiter[0]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[0]));
    MUX21X1 U3258 (.IN1(mask_ff_rr_arbiter[1]), .IN2(next_mask_rr_arbiter[1]), .S(tail_flit_im_output_module[0]), .Q(temp_mask_ff_rr_arbiter[1]));
    MUX21X1 U3259 (.IN1(temp_mask_ff_rr_arbiter), .IN2(1'sb1), .S(arst_value_rr_arbiter), .Q(mask_ff_rr_arbiter[0]));



    BUFX1 U3260 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[0]) );
    BUFX1 U3261 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter11[1]) );
    BUFX1 U3262 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3263 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3264 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    XNOR2X1 U3265 ( .IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter11) );
    MUX21X1 U3266 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U3267 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    INVX1 U3268 ( .A(i_high_prior_arbiter11[0]), .Y(i_0_not_high_prior_arbiter11) );
    MUX21X1 U3269 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter11), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[0]);
    MUX21X1 U3270 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter11[0]), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(raw_grant[1]);
    MUX21X1 U3271 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U3272 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b1), .S(valid_from_im_output_module[7:4][i_high_prior_arbiter11[0]]), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    NAND2X1 U3273 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(_sv2v_jump_high_prior_arbiter11[1]), .QN(nandres_high_prior_arbiter11) );
    MUX21X1 U3274 (.IN1(_sv2v_jump_high_prior_arbiter11[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[0]));
    MUX21X1 U3275 (.IN1(_sv2v_jump_high_prior_arbiter11[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter11), .Q(_sv2v_jump_high_prior_arbiter11[1]));
    HADDX1 U3276 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U3277 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );
    HADDX1 U3278 ( .A0(i_high_prior_arbiter11[0]), .B0(1'b1), .C1(i_high_prior_arbiter11[1]), .SO(i_high_prior_arbiter11[0]) );



    BUFX1 U3279 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[0]) );
    BUFX1 U3280 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter21[1]) );
    BUFX1 U3281 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3282 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3283 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    XNOR2X1 U3284 ( .IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U3285 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U3286 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    INVX1 U3287 ( .A(i_high_prior_arbiter21[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U3288 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[0]);
    MUX21X1 U3289 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter21[0]), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(masked_grant[1]);
    MUX21X1 U3290 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U3291 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter21[0]]), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    NAND2X1 U3292 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(_sv2v_jump_high_prior_arbiter21[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U3293 (.IN1(_sv2v_jump_high_prior_arbiter21[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[0]));
    MUX21X1 U3294 (.IN1(_sv2v_jump_high_prior_arbiter21[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter21[1]));
    HADDX1 U3295 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U3296 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    HADDX1 U3297 ( .A0(i_high_prior_arbiter21[0]), .B0(1'b1), .C1(i_high_prior_arbiter21[1]), .SO(i_high_prior_arbiter21[0]) );
    

    BUFX1 U3298 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[0]) );
    BUFX1 U3299 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter1[1]) );
    AND2X1 U3300 ( .A(mask_ff_rr_arbiter1[0]), .B(valid_from_im_output_module[7:4][0]), .Y(mask_req_rr_arbiter1[0]) );
    AND2X1 U3301 ( .A(mask_ff_rr_arbiter1[1]), .B(valid_from_im_output_module[7:4][1]), .Y(mask_req_rr_arbiter1[1]) );
    BUFX1 U3302 ( .A(mask_ff_rr_arbiter1[0]), .Y(next_mask_rr_arbiter1[0]) );
    BUFX1 U3303 ( .A(mask_ff_rr_arbiter1[1]), .Y(next_mask_rr_arbiter1[1]) );
    XNOR2X1 U3304 ( .IN1(mask_req_rr_arbiter1[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter1) );
    XNOR2X1 U3305 ( .IN1(mask_req_rr_arbiter1[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter1) );
    MUX21X1 U3306 (.IN1(masked_grant_rr_arbiter1[0]), .IN2(raw_grant_rr_arbiter1[0]), .S(xnor0res_rr_arbiter1), .Q(grant_im_output_module[7:4][0]));
    MUX21X1 U3307 (.IN1(masked_grant_rr_arbiter1[1]), .IN2(raw_grant_rr_arbiter1[1]), .S(xnor1res_rr_arbiter1), .Q(grant_im_output_module[7:4][1]));

    BUFX1 U3308 ( .A(1'b0), .Y(i_rr_arbiter1[1]) );
    MUX21X1 U3309 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter1[0]));

    AND2X1 U3310 ( .A(_sv2v_jump_rr_rr_arbiter1[1]), .B(1'b0), .Y(firstif_rr_arbiter1) );
    MUX21X1 U3311 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U3312 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(firstif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    AND2X1 U3313 ( .A(firstif_rr_arbiter1), .B(grant_im_output_module[7:4][i_rr_arbiter1[0]]), .Y(secondif_rr_arbiter1) );
    MUX21X1 U3314 (.IN1(next_mask_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[0]));
    MUX21X1 U3315 (.IN1(next_mask_rr_arbiter1[1]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(next_mask_rr_arbiter1[1]));
    MUX21X1 U3316 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter1[0]), .Q(j_rr_arbiter1[0]));
    AND2X1 U3317 ( .A(secondif_rr_arbiter1), .B(j_rr_arbiter1[0]), .Y(thirdif_rr_arbiter1) );
    MUX21X1 U3318 (.IN1(next_mask_rr_arbiter1[j_rr_arbiter1[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter1), .Q(next_mask_rr_arbiter1[j_rr_arbiter1[0]]));
    MUX21X1 U3319 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U3320 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b1), .S(secondif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));
    NAND2X1 U3321 ( .IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(_sv2v_jump_rr_rr_arbiter1[1]), .QN(fourthif_rr_arbiter1) );
    MUX21X1 U3322 (.IN1(_sv2v_jump_rr_rr_arbiter1[0]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[0]));
    MUX21X1 U3323 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(fourthif_rr_arbiter1), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    MUX21X1 U3324 (.IN1(_sv2v_jump_rr_rr_arbiter1[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter1[1]));

    DFFX2 U3325 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter1) );
    DFFX2 U3326 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter1) );
    MUX21X1 U3327 (.IN1(mask_ff_rr_arbiter1[0]), .IN2(next_mask_rr_arbiter1[0]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[0]));
    MUX21X1 U3328 (.IN1(mask_ff_rr_arbiter1[1]), .IN2(next_mask_rr_arbiter1[1]), .S(tail_flit_im_output_module[1]), .Q(temp_mask_ff_rr_arbiter11[1]));
    MUX21X1 U3329 (.IN1(temp_mask_ff_rr_arbiter11), .IN2(1'sb1), .S(arst_value_rr_arbiter1), .Q(mask_ff_rr_arbiter1[0]));





    BUFX1 U3330 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[0]) );
    BUFX1 U3331 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter12[1]) );
    BUFX1 U3332 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3333 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3334 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    XNOR2X1 U3335 ( .IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter12) );
    MUX21X1 U3336 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U3337 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    INVX1 U3338 ( .A(i_high_prior_arbiter12[0]), .Y(i_0_not_high_prior_arbiter12) );
    MUX21X1 U3339 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter12), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[0]);
    MUX21X1 U3340 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter12[0]), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(raw_grant[1]);
    MUX21X1 U3341 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U3342 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b1), .S(valid_from_im_output_module[11:8][i_high_prior_arbiter12[0]]), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    NAND2X1 U3343 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(_sv2v_jump_high_prior_arbiter12[1]), .QN(nandres_high_prior_arbiter12) );
    MUX21X1 U3344 (.IN1(_sv2v_jump_high_prior_arbiter12[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[0]));
    MUX21X1 U3345 (.IN1(_sv2v_jump_high_prior_arbiter12[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter12), .Q(_sv2v_jump_high_prior_arbiter12[1]));
    HADDX1 U3346 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U3347 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );
    HADDX1 U3348 ( .A0(i_high_prior_arbiter12[0]), .B0(1'b1), .C1(i_high_prior_arbiter12[1]), .SO(i_high_prior_arbiter12[0]) );



    BUFX1 U3349 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[0]) );
    BUFX1 U3350 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter22[1]) );
    BUFX1 U3351 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3352 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3353 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    XNOR2X1 U3354 ( .IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22) );
    MUX21X1 U3355 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U3356 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    INVX1 U3357 ( .A(i_high_prior_arbiter22[0]), .Y(i_0_not_high_prior_arbiter22) );
    MUX21X1 U3358 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[0]);
    MUX21X1 U3359 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter22[0]), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(masked_grant[1]);
    MUX21X1 U3360 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U3361 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter22[0]]), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    NAND2X1 U3362 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(_sv2v_jump_high_prior_arbiter22[1]), .QN(nandres_high_prior_arbiter22) );
    MUX21X1 U3363 (.IN1(_sv2v_jump_high_prior_arbiter22[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[0]));
    MUX21X1 U3364 (.IN1(_sv2v_jump_high_prior_arbiter22[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22), .Q(_sv2v_jump_high_prior_arbiter22[1]));
    HADDX1 U3365 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U3366 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    HADDX1 U3367 ( .A0(i_high_prior_arbiter22[0]), .B0(1'b1), .C1(i_high_prior_arbiter22[1]), .SO(i_high_prior_arbiter22[0]) );
    

    BUFX1 U3368 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[0]) );
    BUFX1 U3369 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter2[1]) );
    AND2X1 U3370 ( .A(mask_ff_rr_arbiter2[0]), .B(valid_from_im_output_module[11:8][0]), .Y(mask_req_rr_arbiter2[0]) );
    AND2X1 U3371 ( .A(mask_ff_rr_arbiter2[1]), .B(valid_from_im_output_module[11:8][1]), .Y(mask_req_rr_arbiter2[1]) );
    BUFX1 U3372 ( .A(mask_ff_rr_arbiter2[0]), .Y(next_mask_rr_arbiter2[0]) );
    BUFX1 U3373 ( .A(mask_ff_rr_arbiter2[1]), .Y(next_mask_rr_arbiter2[1]) );
    XNOR2X1 U3374 ( .IN1(mask_req_rr_arbiter2[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter2) );
    XNOR2X1 U3375 ( .IN1(mask_req_rr_arbiter2[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter2) );
    MUX21X1 U3376 (.IN1(masked_grant_rr_arbiter2[0]), .IN2(raw_grant_rr_arbiter2[0]), .S(xnor0res_rr_arbiter2), .Q(grant_im_output_module[11:8][0]));
    MUX21X1 U3377 (.IN1(masked_grant_rr_arbiter2[1]), .IN2(raw_grant_rr_arbiter2[1]), .S(xnor1res_rr_arbiter2), .Q(grant_im_output_module[11:8][1]));

    BUFX1 U3378 ( .A(1'b0), .Y(i_rr_arbiter2[1]) );
    MUX21X1 U3379 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter2[0]));

    AND2X1 U3380 ( .A(_sv2v_jump_rr_rr_arbiter2[1]), .B(1'b0), .Y(firstif_rr_arbiter2) );
    MUX21X1 U3381 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U3382 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(firstif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    AND2X1 U3383 ( .A(firstif_rr_arbiter2), .B(grant_im_output_module[11:8][i_rr_arbiter2[0]]), .Y(secondif_rr_arbiter2) );
    MUX21X1 U3384 (.IN1(next_mask_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[0]));
    MUX21X1 U3385 (.IN1(next_mask_rr_arbiter2[1]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(next_mask_rr_arbiter2[1]));
    MUX21X1 U3386 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter2[0]), .Q(j_rr_arbiter2[0]));
    AND2X1 U3387 ( .A(secondif_rr_arbiter2), .B(j_rr_arbiter2[0]), .Y(thirdif_rr_arbiter2) );
    MUX21X1 U3388 (.IN1(next_mask_rr_arbiter2[j_rr_arbiter2[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter2), .Q(next_mask_rr_arbiter2[j_rr_arbiter2[0]]));
    MUX21X1 U3389 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U3390 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b1), .S(secondif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));
    NAND2X1 U3391 ( .IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(_sv2v_jump_rr_rr_arbiter2[1]), .QN(fourthif_rr_arbiter2) );
    MUX21X1 U3392 (.IN1(_sv2v_jump_rr_rr_arbiter2[0]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[0]));
    MUX21X1 U3393 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(fourthif_rr_arbiter2), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    MUX21X1 U3394 (.IN1(_sv2v_jump_rr_rr_arbiter2[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter2[1]));

    DFFX2 U3395 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter2) );
    DFFX2 U3396 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter2) );
    MUX21X1 U3397 (.IN1(mask_ff_rr_arbiter2[0]), .IN2(next_mask_rr_arbiter2[0]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[0]));
    MUX21X1 U3398 (.IN1(mask_ff_rr_arbiter2[1]), .IN2(next_mask_rr_arbiter2[1]), .S(tail_flit_im_output_module[2]), .Q(temp_mask_ff_rr_arbiter22[1]));
    MUX21X1 U3399 (.IN1(temp_mask_ff_rr_arbiter22), .IN2(1'sb1), .S(arst_value_rr_arbiter2), .Q(mask_ff_rr_arbiter2[0]));


    XNOR2X1 U3400 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37]), .IN2(vc_channel_output_module[1]), .QN(xnor1resu1_output_module) );
    XNOR2X1 U3401 ( .IN1(int_map_req_v[36:0][in_mod_output_module[1:0]*37-1]), .IN2(vc_channel_output_module[0]), .QN(xnor2resu1_output_module) );
    AND2X1 U3402 ( .IN1(xnor1resu1_output_module), .IN2(xnor2resu1_output_module), .Q(and1resu1_output_module) );
    MUX21X1 U3403 (.IN1(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]), .IN2(1'b1), .S(and1resu1_output_module), .Q(valid_from_im_output_module[(vc_channel_output_module[1:0]*4) + in_mod_output_module[1:0]]);
    HADDX1 U3404 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3405 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3406 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3407 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3408 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3409 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3410 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3411 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3412 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3413 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );  
    HADDX1 U3414 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3415 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3416 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3417 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) ); 
    XOR2X1 U3418 ( .IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .Q(xor1resu1_output_module) );
    MUX21X1 U3419 (.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[0]));
    MUX21X1 U3420 (.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module[1]));
    MUX21X1 U3421 (.IN1(_sv2v_jump_output_module_1[0]), .IN2(_sv2v_jump_output_module[0]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[0]));
    MUX21X1 U3422 (.IN1(_sv2v_jump_output_module_1[1]), .IN2(_sv2v_jump_output_module[1]), .S(xor1resu1_output_module), .Q(_sv2v_jump_output_module_1[1]));
    AND2X1 U3423 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[vc_channel_output_module[1:0]*4+in_mod_output_module[1:0]]), .Q(and2resu1_output_module) );

    MUX21X1 U3424(.IN1(head_flit_output_module[3]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+3]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[3]));
	MUX21X1 U3425(.IN1(head_flit_output_module[4]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+4]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[4]));
	MUX21X1 U3426(.IN1(head_flit_output_module[5]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+5]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[5]));
	MUX21X1 U3427(.IN1(head_flit_output_module[6]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+6]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[6]));
	MUX21X1 U3428(.IN1(head_flit_output_module[7]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+7]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[7]));
	MUX21X1 U3429(.IN1(head_flit_output_module[8]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+8]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[8]));
	MUX21X1 U3430(.IN1(head_flit_output_module[9]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+9]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[9]));
	MUX21X1 U3431(.IN1(head_flit_output_module[10]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+10]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[10]));
	MUX21X1 U3432(.IN1(head_flit_output_module[11]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+11]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[11]));
	MUX21X1 U3433(.IN1(head_flit_output_module[12]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+12]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[12]));
	MUX21X1 U3434(.IN1(head_flit_output_module[13]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+13]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[13]));
	MUX21X1 U3435(.IN1(head_flit_output_module[14]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+14]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[14]));
	MUX21X1 U3436(.IN1(head_flit_output_module[15]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+15]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[15]));
	MUX21X1 U3437(.IN1(head_flit_output_module[16]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+16]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[16]));
	MUX21X1 U3438(.IN1(head_flit_output_module[17]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+17]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[17]));
	MUX21X1 U3439(.IN1(head_flit_output_module[18]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+18]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[18]));
	MUX21X1 U3440(.IN1(head_flit_output_module[19]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+19]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[19]));
	MUX21X1 U3441(.IN1(head_flit_output_module[20]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+20]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[20]));
	MUX21X1 U3442(.IN1(head_flit_output_module[21]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+21]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[21]));
	MUX21X1 U3443(.IN1(head_flit_output_module[22]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+22]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[22]));
	MUX21X1 U3444(.IN1(head_flit_output_module[23]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+23]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[23]));
	MUX21X1 U3445(.IN1(head_flit_output_module[24]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+24]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[24]));
	MUX21X1 U3446(.IN1(head_flit_output_module[25]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+25]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[25]));
	MUX21X1 U3447(.IN1(head_flit_output_module[26]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+26]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[26]));
	MUX21X1 U3448(.IN1(head_flit_output_module[27]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+27]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[27]));
	MUX21X1 U3449(.IN1(head_flit_output_module[28]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+28]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[28]));
	MUX21X1 U3450(.IN1(head_flit_output_module[29]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+29]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[29]));
	MUX21X1 U3451(.IN1(head_flit_output_module[30]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+30]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[30]));
	MUX21X1 U3452(.IN1(head_flit_output_module[31]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+31]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[31]));
	MUX21X1 U3453(.IN1(head_flit_output_module[32]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+32]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[32]));
	MUX21X1 U3454(.IN1(head_flit_output_module[33]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+33]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[33]));
	MUX21X1 U3455(.IN1(head_flit_output_module[34]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+34]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[34]));
	MUX21X1 U3456(.IN1(head_flit_output_module[35]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+35]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[35]));
	MUX21X1 U3457(.IN1(head_flit_output_module[36]), .IN2(int_map_req_v[36:0][in_mod_output_module[1:0]*37+36]), .S(and2resu1_output_module) ,.Q(head_flit_output_module[36]));

    INVX1 U3458 ( .A(head_flit_output_module[32]), .Y(head_flit_output_module_32_not_output_module) );
    AND2X1 U3459 ( .IN1(head_flit_output_module_32_not_output_module), .IN2(head_flit_output_module[33]), .Q(and3resu1_output_module) );
    NOR4X1 U3460 (.IN1(head_flit_output_module[29]), .IN2(head_flit_output_module[28]), .IN3(head_flit_output_module[27]), .IN4(head_flit_output_module[26]), .Q(nor23resu1_output_module) );
    NOR4X1 U3461 (.IN1(head_flit_output_module[25]), .IN2(head_flit_output_module[24]), .IN3(head_flit_output_module[23]), .IN4(head_flit_output_module[22]), .Q(nor23resu2_output_module) );
    AND2X1 U3462 ( .IN1(nor23resu1_output_module), .IN2(nor23resu2_output_module), .Q(and4resu1_output_module) );
    NOR2X1 U3463 (.IN1(head_flit_output_module[33]), .IN2(head_flit_output_module[32]), .Q(nor23resu3_output_module) );
    AND2X1 U3464 ( .IN1(nor23resu3_output_module), .IN2(and4resu1_output_module), .Q(and5resu1_output_module) );    
    OR2X1 U3465 (.IN1(and3resu1_output_module), .IN2(nor23resu3_output_module), .Q(or12resu12_output_module) );
    AND2X1 U3466 ( .IN1(ext_resp_v_i[1:0][0]), .IN2(or12resu12_output_module), .Q(and6resu1_output_module) );    
	MUX21X1 U3467(.IN1(tail_flit_im_output_module[vc_channel_output_module[1:0]]), .IN2(and6resu1_output_module), .S(and2resu1_output_module) ,.Q(tail_flit_im_output_module[vc_channel_output_module[1:0]]);
	MUX21X1 U3468(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3469(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and2resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
    NAND2X1 U3470(.A(_sv2v_jump_output_module[0]),.B(_sv2v_jump_output_module[1]),.Y(nand1resu_output_module));

    AND2X1 U3471 ( .IN1(xor1resu1_output_module), .IN2(nand1resu_output_module), .Q(and7resu1) );    
	MUX21X1 U3472(.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3473(.IN1(_sv2v_jump_output_module[1]), .IN2(_sv2v_jump_output_module_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	MUX21X1 U3474(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3475(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module[1]);

	HADDX1 U3476 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3477 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3478 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3479 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3480 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U3481 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3482 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3483 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3484 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3485 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
	HADDX1 U3486 ( .A0(vc_channel_output_module[0]), .B0(1'b1), .C1(vc_channel_output_module[1]), .SO(vc_channel_output_module[0]) );
    HADDX1 U3487 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3488 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3489 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );
    HADDX1 U3490 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(in_mod_output_module[1]), .SO(in_mod_output_module[0]) );



	BUFX1 U3491(.A(1'b0), .Y(_sv2v_jump_output_module[0]));
	BUFX1 U3492(.A(1'b0), .Y(_sv2v_jump_output_module[1]));
    AND2X1 U3493 ( .IN1(xor1resu1_output_module), .IN2(grant_im_output_module[i_output_module[1:0] * 4+:4]), .Q(and8resu1_output_module) );    
    MUX21X1 U3494(.IN1(vc_ch_act_out_output_module[0]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[0]);
	MUX21X1 U3495(.IN1(vc_ch_act_out_output_module[1]), .IN2(i_output_module[1:0]), .S(and8resu1_output_module) ,.Q(vc_ch_act_out_output_module[1]);
	MUX21X1 U3496(.IN1(req_out_output_module), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(req_out_output_module);
	MUX21X1 U3497(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3498(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and8resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);
	HADDX1 U3499 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U3500 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    HADDX1 U3501 ( .A0(in_mod_output_module[0]), .B0(1'b1), .C1(i_output_module[1]), .SO(i_output_module[0]) );

    NOR2X1 U3502 (.IN1(_sv2v_jump_output_module[0]), .IN2(_sv2v_jump_output_module[1]), .Q(norfinresu1_output_module) );
    AND2X1 U3503 ( .IN1(norfinresu1_output_module), .IN2(req_out_output_module), .Q(and9resu1_output_module) );    
	HADDX1 U3504 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module[1]), .SO(i_output_module[0]) );
    AND2X1 U3505 ( .IN1(and9resu1_output_module), .IN2(grant_im_output_module[(vc_ch_act_out_output_module * 4) + i_output_module[1:0]]), .Q(and10resu1_output_module) );    

	MUX21X1 U3506(.IN1(ext_req_v_o[36:0][3]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+3]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][3]));
	MUX21X1 U3507(.IN1(ext_req_v_o[36:0][4]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+4]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][4]));
	MUX21X1 U3508(.IN1(ext_req_v_o[36:0][5]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+5]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][5]));
	MUX21X1 U3509(.IN1(ext_req_v_o[36:0][6]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+6]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][6]));
	MUX21X1 U3510(.IN1(ext_req_v_o[36:0][7]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+7]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][7]));
	MUX21X1 U3511(.IN1(ext_req_v_o[36:0][8]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+8]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][8]));
	MUX21X1 U3512(.IN1(ext_req_v_o[36:0][9]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+9]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][9]));
	MUX21X1 U3513(.IN1(ext_req_v_o[36:0][10]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+10]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][10]));
	MUX21X1 U3514(.IN1(ext_req_v_o[36:0][11]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+11]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][11]));
	MUX21X1 U3515(.IN1(ext_req_v_o[36:0][12]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+12]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][12]));
	MUX21X1 U3516(.IN1(ext_req_v_o[36:0][13]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+13]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][13]));
	MUX21X1 U3517(.IN1(ext_req_v_o[36:0][14]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+14]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][14]));
	MUX21X1 U3518(.IN1(ext_req_v_o[36:0][15]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+15]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][15]));
	MUX21X1 U3519(.IN1(ext_req_v_o[36:0][16]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+16]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][16]));
	MUX21X1 U3520(.IN1(ext_req_v_o[36:0][17]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+17]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][17]));
	MUX21X1 U3521(.IN1(ext_req_v_o[36:0][18]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+18]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][18]));
	MUX21X1 U3522(.IN1(ext_req_v_o[36:0][19]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+19]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][19]));
	MUX21X1 U3523(.IN1(ext_req_v_o[36:0][20]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+20]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][20]));
	MUX21X1 U3524(.IN1(ext_req_v_o[36:0][21]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+21]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][21]));
	MUX21X1 U3525(.IN1(ext_req_v_o[36:0][22]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+22]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][22]));
	MUX21X1 U3526(.IN1(ext_req_v_o[36:0][23]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+23]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][23]));
	MUX21X1 U3527(.IN1(ext_req_v_o[36:0][24]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+24]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][24]));
	MUX21X1 U3528(.IN1(ext_req_v_o[36:0][25]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+25]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][25]));
	MUX21X1 U3529(.IN1(ext_req_v_o[36:0][26]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+26]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][26]));
	MUX21X1 U3530(.IN1(ext_req_v_o[36:0][27]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+27]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][27]));
	MUX21X1 U3531(.IN1(ext_req_v_o[36:0][28]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+28]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][28]));
	MUX21X1 U3532(.IN1(ext_req_v_o[36:0][29]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+29]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][29]));
	MUX21X1 U3533(.IN1(ext_req_v_o[36:0][30]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+30]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][30]));
	MUX21X1 U3534(.IN1(ext_req_v_o[36:0][31]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+31]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][31]));
	MUX21X1 U3535(.IN1(ext_req_v_o[36:0][32]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+32]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][32]));
	MUX21X1 U3536(.IN1(ext_req_v_o[36:0][33]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+33]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][33]));
	MUX21X1 U3537(.IN1(ext_req_v_o[36:0][34]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+34]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][34]));
	MUX21X1 U3538(.IN1(ext_req_v_o[36:0][35]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+35]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][35]));
	MUX21X1 U3539(.IN1(ext_req_v_o[36:0][36]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37+36]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][36]));

	MUX21X1 U3540(.IN1(ext_req_v_o[36:0][0]), .IN2(int_map_req_v[36:0][i_output_module[1:0]*37]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][0]);
	MUX21X1 U3541(.IN1(ext_req_v_o[36:0][1]), .IN2(vc_ch_act_out_output_module[0]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][1]);
	MUX21X1 U3542(.IN1(ext_req_v_o[36:0][2]), .IN2(vc_ch_act_out_output_module[1]), .S(and10resu1_output_module) ,.Q(ext_req_v_o[36:0][2]);    
	MUX21X1 U3543(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3544(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b1), .S(and10resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);    

    AND2X1 U3545 ( .IN1(and9resu1_output_module), .IN2(nand1resu_output_module), .Q(and11resu1_output_module) );    
	MUX21X1 U3546(.IN1(_sv2v_jump_output_module[0]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[0]);
	MUX21X1 U3547(.IN1(_sv2v_jump_output_module[1]), .IN2(1'b0), .S(and11resu1_output_module) ,.Q(_sv2v_jump_output_module[1]);  





    BUFX1 U3548 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[0]) );
    BUFX1 U3549 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter111[1]) );
    BUFX1 U3550 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3551 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3552 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    XNOR2X1 U3553 ( .IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter111) );
    MUX21X1 U3554 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U3555 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    INVX1 U3556 ( .A(i_high_prior_arbiter111[0]), .Y(i_0_not_high_prior_arbiter111) );
    MUX21X1 U3557 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter111), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[0]);
    MUX21X1 U3558 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter111[0]), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(raw_grant[1]);
    MUX21X1 U3559 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U3560 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[3:0][i_high_prior_arbiter111[0]]), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    NAND2X1 U3561 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(_sv2v_jump_high_prior_arbiter111[1]), .QN(nandres_high_prior_arbiter111) );
    MUX21X1 U3562 (.IN1(_sv2v_jump_high_prior_arbiter111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[0]));
    MUX21X1 U3563 (.IN1(_sv2v_jump_high_prior_arbiter111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter111), .Q(_sv2v_jump_high_prior_arbiter111[1]));
    HADDX1 U3564 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U3565 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );
    HADDX1 U3566 ( .A0(i_high_prior_arbiter111[0]), .B0(1'b1), .C1(i_high_prior_arbiter111[1]), .SO(i_high_prior_arbiter111[0]) );



    BUFX1 U3567 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[0]) );
    BUFX1 U3568 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter211[1]) );
    BUFX1 U3569 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3570 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3571 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    XNOR2X1 U3572 ( .IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter21) );
    MUX21X1 U3573 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U3574 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    INVX1 U3575 ( .A(i_high_prior_arbiter211[0]), .Y(i_0_not_high_prior_arbiter21) );
    MUX21X1 U3576 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter21), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[0]);
    MUX21X1 U3577 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter211[0]), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(masked_grant[1]);
    MUX21X1 U3578 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U3579 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter211[0]]), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    NAND2X1 U3580 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(_sv2v_jump_high_prior_arbiter211[1]), .QN(nandres_high_prior_arbiter21) );
    MUX21X1 U3581 (.IN1(_sv2v_jump_high_prior_arbiter211[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[0]));
    MUX21X1 U3582 (.IN1(_sv2v_jump_high_prior_arbiter211[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter21), .Q(_sv2v_jump_high_prior_arbiter211[1]));
    HADDX1 U3583 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U3584 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    HADDX1 U3585 ( .A0(i_high_prior_arbiter211[0]), .B0(1'b1), .C1(i_high_prior_arbiter211[1]), .SO(i_high_prior_arbiter211[0]) );
    

    BUFX1 U3586 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[0]) );
    BUFX1 U3587 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter11[1]) );
    AND2X1 U3588 ( .A(mask_ff_rr_arbiter11[0]), .B(valid_from_im_output_module1[3:0][0]), .Y(mask_req_rr_arbiter11[0]) );
    AND2X1 U3589 ( .A(mask_ff_rr_arbiter11[1]), .B(valid_from_im_output_module1[3:0][1]), .Y(mask_req_rr_arbiter11[1]) );
    BUFX1 U3590 ( .A(mask_ff_rr_arbiter11[0]), .Y(next_mask_rr_arbiter11[0]) );
    BUFX1 U3591 ( .A(mask_ff_rr_arbiter11[1]), .Y(next_mask_rr_arbiter11[1]) );
    XNOR2X1 U3592 ( .IN1(mask_req_rr_arbiter11[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter11) );
    XNOR2X1 U3593 ( .IN1(mask_req_rr_arbiter11[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter11) );
    MUX21X1 U3594 (.IN1(masked_grant_rr_arbiter11[0]), .IN2(raw_grant_rr_arbiter11[0]), .S(xnor0res_rr_arbiter11), .Q(grant_im_output_module1[3:0][0]));
    MUX21X1 U3595 (.IN1(masked_grant_rr_arbiter11[1]), .IN2(raw_grant_rr_arbiter11[1]), .S(xnor1res_rr_arbiter11), .Q(grant_im_output_module1[3:0][1]));

    BUFX1 U3596 ( .A(1'b0), .Y(i_rr_arbiter11[1]) );
    MUX21X1 U3597 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter11[0]));

    AND2X1 U3598 ( .A(_sv2v_jump_rr_rr_arbiter11[1]), .B(1'b0), .Y(firstif_rr_arbiter11) );
    MUX21X1 U3599 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U3600 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(firstif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    AND2X1 U3601 ( .A(firstif_rr_arbiter11), .B(grant_im_output_module1[3:0][i_rr_arbiter11[0]]), .Y(secondif_rr_arbiter11) );
    MUX21X1 U3602 (.IN1(next_mask_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[0]));
    MUX21X1 U3603 (.IN1(next_mask_rr_arbiter11[1]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(next_mask_rr_arbiter11[1]));
    MUX21X1 U3604 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter11[0]), .Q(j_rr_arbiter11[0]));
    AND2X1 U3605 ( .A(secondif_rr_arbiter11), .B(j_rr_arbiter11[0]), .Y(thirdif_rr_arbiter11) );
    MUX21X1 U3606 (.IN1(next_mask_rr_arbiter11[j_rr_arbiter11[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter11), .Q(next_mask_rr_arbiter11[j_rr_arbiter11[0]]));
    MUX21X1 U3607 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U3608 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b1), .S(secondif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));
    NAND2X1 U3609 ( .IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(_sv2v_jump_rr_rr_arbiter11[1]), .QN(fourthif_rr_arbiter11) );
    MUX21X1 U3610 (.IN1(_sv2v_jump_rr_rr_arbiter11[0]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[0]));
    MUX21X1 U3611 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(fourthif_rr_arbiter11), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    MUX21X1 U3612 (.IN1(_sv2v_jump_rr_rr_arbiter11[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter11[1]));

    DFFX2 U3613 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter11) );
    DFFX2 U3614 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter11) );
    MUX21X1 U3615 (.IN1(mask_ff_rr_arbiter11[0]), .IN2(next_mask_rr_arbiter11[0]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[0]));
    MUX21X1 U3616 (.IN1(mask_ff_rr_arbiter11[1]), .IN2(next_mask_rr_arbiter11[1]), .S(tail_flit_im_output_module1[0]), .Q(temp_mask_ff_rr_arbiter1111[1]));
    MUX21X1 U3617 (.IN1(temp_mask_ff_rr_arbiter1111), .IN2(1'sb1), .S(arst_value_rr_arbiter11), .Q(mask_ff_rr_arbiter11[0]));



    BUFX1 U3618 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[0]) );
    BUFX1 U3619 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1111[1]) );
    BUFX1 U3620 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3621 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3622 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    XNOR2X1 U3623 ( .IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1111) );
    MUX21X1 U3624 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U3625 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    INVX1 U3626 ( .A(i_high_prior_arbiter1111[0]), .Y(i_0_not_high_prior_arbiter1111) );
    MUX21X1 U3627 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1111), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[0]);
    MUX21X1 U3628 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1111[0]), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(raw_grant[1]);
    MUX21X1 U3629 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U3630 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b1), .S(valid_from_im_output_module1[7:4][i_high_prior_arbiter1111[0]]), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    NAND2X1 U3631 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(_sv2v_jump_high_prior_arbiter1111[1]), .QN(nandres_high_prior_arbiter1111) );
    MUX21X1 U3632 (.IN1(_sv2v_jump_high_prior_arbiter1111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[0]));
    MUX21X1 U3633 (.IN1(_sv2v_jump_high_prior_arbiter1111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1111), .Q(_sv2v_jump_high_prior_arbiter1111[1]));
    HADDX1 U3634 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U3635 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );
    HADDX1 U3636 ( .A0(i_high_prior_arbiter1111[0]), .B0(1'b1), .C1(i_high_prior_arbiter1111[1]), .SO(i_high_prior_arbiter1111[0]) );



    BUFX1 U3637 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[0]) );
    BUFX1 U3638 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2111[1]) );
    BUFX1 U3639 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3640 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3641 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    XNOR2X1 U3642 ( .IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2111) );
    MUX21X1 U3643 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U3644 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    INVX1 U3645 ( .A(i_high_prior_arbiter2111[0]), .Y(i_0_not_high_prior_arbiter2111) );
    MUX21X1 U3646 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2111), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[0]);
    MUX21X1 U3647 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2111[0]), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(masked_grant[1]);
    MUX21X1 U3648 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U3649 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2111[0]]), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    NAND2X1 U3650 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(_sv2v_jump_high_prior_arbiter2111[1]), .QN(nandres_high_prior_arbiter2111) );
    MUX21X1 U3651 (.IN1(_sv2v_jump_high_prior_arbiter2111[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[0]));
    MUX21X1 U3652 (.IN1(_sv2v_jump_high_prior_arbiter2111[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2111), .Q(_sv2v_jump_high_prior_arbiter2111[1]));
    HADDX1 U3653 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U3654 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    HADDX1 U3655 ( .A0(i_high_prior_arbiter2111[0]), .B0(1'b1), .C1(i_high_prior_arbiter2111[1]), .SO(i_high_prior_arbiter2111[0]) );
    

    BUFX1 U3656 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[0]) );
    BUFX1 U3657 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter111[1]) );
    AND2X1 U3658 ( .A(mask_ff_rr_arbiter111[0]), .B(valid_from_im_output_module1[7:4][0]), .Y(mask_req_rr_arbiter111[0]) );
    AND2X1 U3659 ( .A(mask_ff_rr_arbiter111[1]), .B(valid_from_im_output_module1[7:4][1]), .Y(mask_req_rr_arbiter111[1]) );
    BUFX1 U3660 ( .A(mask_ff_rr_arbiter111[0]), .Y(next_mask_rr_arbiter111[0]) );
    BUFX1 U3661 ( .A(mask_ff_rr_arbiter111[1]), .Y(next_mask_rr_arbiter111[1]) );
    XNOR2X1 U3662 ( .IN1(mask_req_rr_arbiter111[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter111) );
    XNOR2X1 U3663 ( .IN1(mask_req_rr_arbiter111[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter111) );
    MUX21X1 U3664 (.IN1(masked_grant_rr_arbiter111[0]), .IN2(raw_grant_rr_arbiter111[0]), .S(xnor0res_rr_arbiter111), .Q(grant_im_output_module1[7:4][0]));
    MUX21X1 U3665 (.IN1(masked_grant_rr_arbiter111[1]), .IN2(raw_grant_rr_arbiter111[1]), .S(xnor1res_rr_arbiter111), .Q(grant_im_output_module1[7:4][1]));

    BUFX1 U3666 ( .A(1'b0), .Y(i_rr_arbiter111[1]) );
    MUX21X1 U3667 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter111[0]));

    AND2X1 U3668 ( .A(_sv2v_jump_rr_rr_arbiter111[1]), .B(1'b0), .Y(firstif_rr_arbiter111) );
    MUX21X1 U3669 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U3670 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(firstif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    AND2X1 U3671 ( .A(firstif_rr_arbiter111), .B(grant_im_output_module1[7:4][i_rr_arbiter111[0]]), .Y(secondif_rr_arbiter111) );
    MUX21X1 U3672 (.IN1(next_mask_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[0]));
    MUX21X1 U3673 (.IN1(next_mask_rr_arbiter111[1]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(next_mask_rr_arbiter111[1]));
    MUX21X1 U3674 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter111[0]), .Q(j_rr_arbiter111[0]));
    AND2X1 U3675 ( .A(secondif_rr_arbiter111), .B(j_rr_arbiter111[0]), .Y(thirdif_rr_arbiter111) );
    MUX21X1 U3676 (.IN1(next_mask_rr_arbiter111[j_rr_arbiter111[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter111), .Q(next_mask_rr_arbiter111[j_rr_arbiter111[0]]));
    MUX21X1 U3677 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U3678 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b1), .S(secondif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));
    NAND2X1 U3679 ( .IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(_sv2v_jump_rr_rr_arbiter111[1]), .QN(fourthif_rr_arbiter111) );
    MUX21X1 U3680 (.IN1(_sv2v_jump_rr_rr_arbiter111[0]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[0]));
    MUX21X1 U3681 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(fourthif_rr_arbiter111), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    MUX21X1 U3682 (.IN1(_sv2v_jump_rr_rr_arbiter111[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter111[1]));

    DFFX2 U3683 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter111) );
    DFFX2 U3684 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter111) );
    MUX21X1 U3685 (.IN1(mask_ff_rr_arbiter111[0]), .IN2(next_mask_rr_arbiter111[0]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[0]));
    MUX21X1 U3686 (.IN1(mask_ff_rr_arbiter111[1]), .IN2(next_mask_rr_arbiter111[1]), .S(tail_flit_im_output_module1[1]), .Q(temp_mask_ff_rr_arbiter111111[1]));
    MUX21X1 U3687 (.IN1(temp_mask_ff_rr_arbiter111111), .IN2(1'sb1), .S(arst_value_rr_arbiter111), .Q(mask_ff_rr_arbiter111[0]));





    BUFX1 U3688 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[0]) );
    BUFX1 U3689 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1112[1]) );
    BUFX1 U3690 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3691 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3692 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    XNOR2X1 U3693 ( .IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1112) );
    MUX21X1 U3694 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U3695 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    INVX1 U3696 ( .A(i_high_prior_arbiter1112[0]), .Y(i_0_not_high_prior_arbiter1112) );
    MUX21X1 U3697 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1112), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[0]);
    MUX21X1 U3698 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1112[0]), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(raw_grant[1]);
    MUX21X1 U3699 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U3700 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b1), .S(valid_from_im_output_module1[11:8][i_high_prior_arbiter1112[0]]), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    NAND2X1 U3701 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(_sv2v_jump_high_prior_arbiter1112[1]), .QN(nandres_high_prior_arbiter1112) );
    MUX21X1 U3702 (.IN1(_sv2v_jump_high_prior_arbiter1112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[0]));
    MUX21X1 U3703 (.IN1(_sv2v_jump_high_prior_arbiter1112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1112), .Q(_sv2v_jump_high_prior_arbiter1112[1]));
    HADDX1 U3704 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U3705 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );
    HADDX1 U3706 ( .A0(i_high_prior_arbiter1112[0]), .B0(1'b1), .C1(i_high_prior_arbiter1112[1]), .SO(i_high_prior_arbiter1112[0]) );



    BUFX1 U3707 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[0]) );
    BUFX1 U3708 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2112[1]) );
    BUFX1 U3709 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3710 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3711 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    XNOR2X1 U3712 ( .IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter212) );
    MUX21X1 U3713 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U3714 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    INVX1 U3715 ( .A(i_high_prior_arbiter2112[0]), .Y(i_0_not_high_prior_arbiter212) );
    MUX21X1 U3716 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter212), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[0]);
    MUX21X1 U3717 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2112[0]), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(masked_grant[1]);
    MUX21X1 U3718 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U3719 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2112[0]]), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    NAND2X1 U3720 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(_sv2v_jump_high_prior_arbiter2112[1]), .QN(nandres_high_prior_arbiter212) );
    MUX21X1 U3721 (.IN1(_sv2v_jump_high_prior_arbiter2112[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[0]));
    MUX21X1 U3722 (.IN1(_sv2v_jump_high_prior_arbiter2112[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter212), .Q(_sv2v_jump_high_prior_arbiter2112[1]));
    HADDX1 U3723 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U3724 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    HADDX1 U3725 ( .A0(i_high_prior_arbiter2112[0]), .B0(1'b1), .C1(i_high_prior_arbiter2112[1]), .SO(i_high_prior_arbiter2112[0]) );
    

    BUFX1 U3726 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[0]) );
    BUFX1 U3727 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter112[1]) );
    AND2X1 U3728 ( .A(mask_ff_rr_arbiter112[0]), .B(valid_from_im_output_module1[11:8][0]), .Y(mask_req_rr_arbiter112[0]) );
    AND2X1 U3729 ( .A(mask_ff_rr_arbiter112[1]), .B(valid_from_im_output_module1[11:8][1]), .Y(mask_req_rr_arbiter112[1]) );
    BUFX1 U3730 ( .A(mask_ff_rr_arbiter112[0]), .Y(next_mask_rr_arbiter112[0]) );
    BUFX1 U3731 ( .A(mask_ff_rr_arbiter112[1]), .Y(next_mask_rr_arbiter112[1]) );
    XNOR2X1 U3732 ( .IN1(mask_req_rr_arbiter112[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter112) );
    XNOR2X1 U3733 ( .IN1(mask_req_rr_arbiter112[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter112) );
    MUX21X1 U3734 (.IN1(masked_grant_rr_arbiter112[0]), .IN2(raw_grant_rr_arbiter112[0]), .S(xnor0res_rr_arbiter112), .Q(grant_im_output_module1[11:8][0]));
    MUX21X1 U3735 (.IN1(masked_grant_rr_arbiter112[1]), .IN2(raw_grant_rr_arbiter112[1]), .S(xnor1res_rr_arbiter112), .Q(grant_im_output_module1[11:8][1]));

    BUFX1 U3736 ( .A(1'b0), .Y(i_rr_arbiter112[1]) );
    MUX21X1 U3737 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter112[0]));

    AND2X1 U3738 ( .A(_sv2v_jump_rr_rr_arbiter112[1]), .B(1'b0), .Y(firstif_rr_arbiter112) );
    MUX21X1 U3739 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U3740 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(firstif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    AND2X1 U3741 ( .A(firstif_rr_arbiter112), .B(grant_im_output_module1[11:8][i_rr_arbiter112[0]]), .Y(secondif_rr_arbiter112) );
    MUX21X1 U3742 (.IN1(next_mask_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[0]));
    MUX21X1 U3743 (.IN1(next_mask_rr_arbiter112[1]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(next_mask_rr_arbiter112[1]));
    MUX21X1 U3744 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter112[0]), .Q(j_rr_arbiter112[0]));
    AND2X1 U3745 ( .A(secondif_rr_arbiter112), .B(j_rr_arbiter112[0]), .Y(thirdif_rr_arbiter112) );
    MUX21X1 U3746 (.IN1(next_mask_rr_arbiter112[j_rr_arbiter112[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter112), .Q(next_mask_rr_arbiter112[j_rr_arbiter112[0]]));
    MUX21X1 U3747 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U3748 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b1), .S(secondif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));
    NAND2X1 U3749 ( .IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(_sv2v_jump_rr_rr_arbiter112[1]), .QN(fourthif_rr_arbiter112) );
    MUX21X1 U3750 (.IN1(_sv2v_jump_rr_rr_arbiter112[0]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[0]));
    MUX21X1 U3751 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(fourthif_rr_arbiter112), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    MUX21X1 U3752 (.IN1(_sv2v_jump_rr_rr_arbiter112[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter112[1]));

    DFFX2 U3753 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter112) );
    DFFX2 U3754 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter112) );
    MUX21X1 U3755 (.IN1(mask_ff_rr_arbiter112[0]), .IN2(next_mask_rr_arbiter112[0]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[0]));
    MUX21X1 U3756 (.IN1(mask_ff_rr_arbiter112[1]), .IN2(next_mask_rr_arbiter112[1]), .S(tail_flit_im_output_module1[2]), .Q(temp_mask_ff_rr_arbiter111122[1]));
    MUX21X1 U3757 (.IN1(temp_mask_ff_rr_arbiter111122), .IN2(1'sb1), .S(arst_value_rr_arbiter112), .Q(mask_ff_rr_arbiter112[0]));


    XNOR2X1 U3758 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37]), .IN2(vc_channel_output_module1[1]), .QN(xnor1resu1_output_module1) );
    XNOR2X1 U3759 ( .IN1(int_map_req_v[184:148][in_mod_output_module1[1:0]*37-1]), .IN2(vc_channel_output_module1[0]), .QN(xnor2resu1_output_module1) );
    AND2X1 U3760 ( .IN1(xnor1resu1_output_module1), .IN2(xnor2resu1_output_module1), .Q(and1resu1_output_module1) );
    MUX21X1 U3761 (.IN1(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]), .IN2(1'b1), .S(and1resu1_output_module1), .Q(valid_from_im_output_module1[(vc_channel_output_module1[1:0]*4) + in_mod_output_module1[1:0]]);
    HADDX1 U3762 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3763 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3764 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3765 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3766 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3767 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3768 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3769 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3770 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3771 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );  
    HADDX1 U3772 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3773 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3774 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3775 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) ); 
    XOR2X1 U3776 ( .IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .Q(xor1resu1_output_module1) );
    MUX21X1 U3777 (.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[0]));
    MUX21X1 U3778 (.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1[1]));
    MUX21X1 U3779 (.IN1(_sv2v_jump_output_module1_1[0]), .IN2(_sv2v_jump_output_module1[0]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[0]));
    MUX21X1 U3780 (.IN1(_sv2v_jump_output_module1_1[1]), .IN2(_sv2v_jump_output_module1[1]), .S(xor1resu1_output_module1), .Q(_sv2v_jump_output_module1_1[1]));
    AND2X1 U3781 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[vc_channel_output_module1[1:0]*4+in_mod_output_module1[1:0]]), .Q(and2resu1_output_module1) );

    MUX21X1 U3782(.IN1(head_flit_output_module1[3]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+3]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[3]));
    MUX21X1 U3783(.IN1(head_flit_output_module1[4]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+4]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[4]));
    MUX21X1 U3784(.IN1(head_flit_output_module1[5]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+5]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[5]));
    MUX21X1 U3785(.IN1(head_flit_output_module1[6]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+6]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[6]));
    MUX21X1 U3786(.IN1(head_flit_output_module1[7]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+7]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[7]));
    MUX21X1 U3787(.IN1(head_flit_output_module1[8]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+8]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[8]));
    MUX21X1 U3788(.IN1(head_flit_output_module1[9]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+9]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[9]));
    MUX21X1 U3789(.IN1(head_flit_output_module1[10]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+10]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[10]));
    MUX21X1 U3790(.IN1(head_flit_output_module1[11]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+11]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[11]));
    MUX21X1 U3791(.IN1(head_flit_output_module1[12]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+12]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[12]));
    MUX21X1 U3792(.IN1(head_flit_output_module1[13]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+13]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[13]));
    MUX21X1 U3793(.IN1(head_flit_output_module1[14]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+14]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[14]));
    MUX21X1 U3794(.IN1(head_flit_output_module1[15]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+15]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[15]));
    MUX21X1 U3795(.IN1(head_flit_output_module1[16]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+16]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[16]));
    MUX21X1 U3796(.IN1(head_flit_output_module1[17]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+17]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[17]));
    MUX21X1 U3797(.IN1(head_flit_output_module1[18]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+18]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[18]));
    MUX21X1 U3798(.IN1(head_flit_output_module1[19]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+19]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[19]));
    MUX21X1 U3799(.IN1(head_flit_output_module1[20]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+20]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[20]));
    MUX21X1 U3800(.IN1(head_flit_output_module1[21]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+21]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[21]));
    MUX21X1 U3801(.IN1(head_flit_output_module1[22]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+22]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[22]));
    MUX21X1 U3802(.IN1(head_flit_output_module1[23]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+23]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[23]));
    MUX21X1 U3803(.IN1(head_flit_output_module1[24]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+24]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[24]));
    MUX21X1 U3804(.IN1(head_flit_output_module1[25]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+25]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[25]));
    MUX21X1 U3805(.IN1(head_flit_output_module1[26]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+26]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[26]));
    MUX21X1 U3806(.IN1(head_flit_output_module1[27]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+27]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[27]));
    MUX21X1 U3807(.IN1(head_flit_output_module1[28]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+28]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[28]));
    MUX21X1 U3808(.IN1(head_flit_output_module1[29]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+29]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[29]));
    MUX21X1 U3809(.IN1(head_flit_output_module1[30]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+30]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[30]));
    MUX21X1 U3810(.IN1(head_flit_output_module1[31]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+31]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[31]));
    MUX21X1 U3811(.IN1(head_flit_output_module1[32]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+32]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[32]));
    MUX21X1 U3812(.IN1(head_flit_output_module1[33]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+33]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[33]));
    MUX21X1 U3813(.IN1(head_flit_output_module1[34]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+34]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[34]));
    MUX21X1 U3814(.IN1(head_flit_output_module1[35]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+35]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[35]));
    MUX21X1 U3815(.IN1(head_flit_output_module1[36]), .IN2(int_map_req_v[184:148][in_mod_output_module1[1:0]*37+36]), .S(and2resu1_output_module1) ,.Q(head_flit_output_module1[36]));

    INVX1 U3816 ( .A(head_flit_output_module1[32]), .Y(head_flit_output_module1_32_not_output_module1) );
    AND2X1 U3817 ( .IN1(head_flit_output_module1_32_not_output_module1), .IN2(head_flit_output_module1[33]), .Q(and3resu1_output_module1) );
    NOR4X1 U3818 (.IN1(head_flit_output_module1[29]), .IN2(head_flit_output_module1[28]), .IN3(head_flit_output_module1[27]), .IN4(head_flit_output_module1[26]), .Q(nor23resu1_output_module1) );
    NOR4X1 U3819 (.IN1(head_flit_output_module1[25]), .IN2(head_flit_output_module1[24]), .IN3(head_flit_output_module1[23]), .IN4(head_flit_output_module1[22]), .Q(nor23resu2_output_module1) );
    AND2X1 U3820 ( .IN1(nor23resu1_output_module1), .IN2(nor23resu2_output_module1), .Q(and4resu1_output_module1) );
    NOR2X1 U3821 (.IN1(head_flit_output_module1[33]), .IN2(head_flit_output_module1[32]), .Q(nor23resu3_output_module1) );
    AND2X1 U3822 ( .IN1(nor23resu3_output_module1), .IN2(and4resu1_output_module1), .Q(and5resu1_output_module1) );    
    OR2X1 U3823 (.IN1(and3resu1_output_module1), .IN2(nor23resu3_output_module1), .Q(or12resu12_output_module1) );
    AND2X1 U3824 ( .IN1(ext_resp_v_i[2:1][0]), .IN2(or12resu12_output_module1), .Q(and6resu1_output_module1) );    
    MUX21X1 U3825(.IN1(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]), .IN2(and6resu1_output_module1), .S(and2resu1_output_module1) ,.Q(tail_flit_im_output_module1[vc_channel_output_module1[1:0]]);
    MUX21X1 U3826(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3827(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and2resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    NAND2X1 U3828(.A(_sv2v_jump_output_module1[0]),.B(_sv2v_jump_output_module1[1]),.Y(nand1resu_output_module1));

    AND2X1 U3829 ( .IN1(xor1resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and7resu1) );    
    MUX21X1 U3830(.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3831(.IN1(_sv2v_jump_output_module1[1]), .IN2(_sv2v_jump_output_module1_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    MUX21X1 U3832(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3833(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module1[1]);

    HADDX1 U3834 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3835 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3836 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3837 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3838 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3839 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3840 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3841 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3842 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3843 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3844 ( .A0(vc_channel_output_module1[0]), .B0(1'b1), .C1(vc_channel_output_module1[1]), .SO(vc_channel_output_module1[0]) );
    HADDX1 U3845 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3846 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3847 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );
    HADDX1 U3848 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(in_mod_output_module1[1]), .SO(in_mod_output_module1[0]) );



    BUFX1 U3849(.A(1'b0), .Y(_sv2v_jump_output_module1[0]));
    BUFX1 U3850(.A(1'b0), .Y(_sv2v_jump_output_module1[1]));
    AND2X1 U3851 ( .IN1(xor1resu1_output_module1), .IN2(grant_im_output_module1[i_output_module1[1:0] * 4+:4]), .Q(and8resu1_output_module1) );    
    MUX21X1 U3852(.IN1(vc_ch_act_out_output_module1[0]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[0]);
    MUX21X1 U3853(.IN1(vc_ch_act_out_output_module1[1]), .IN2(i_output_module1[1:0]), .S(and8resu1_output_module1) ,.Q(vc_ch_act_out_output_module1[1]);
    MUX21X1 U3854(.IN1(req_out_output_module1), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(req_out_output_module1);
    MUX21X1 U3855(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3856(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and8resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);
    HADDX1 U3857 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U3858 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    HADDX1 U3859 ( .A0(in_mod_output_module1[0]), .B0(1'b1), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );

    NOR2X1 U3860 (.IN1(_sv2v_jump_output_module1[0]), .IN2(_sv2v_jump_output_module1[1]), .Q(norfinresu1_output_module1) );
    AND2X1 U3861 ( .IN1(norfinresu1_output_module1), .IN2(req_out_output_module1), .Q(and9resu1_output_module1) );    
    HADDX1 U3862 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module1[1]), .SO(i_output_module1[0]) );
    AND2X1 U3863 ( .IN1(and9resu1_output_module1), .IN2(grant_im_output_module1[(vc_ch_act_out_output_module1 * 4) + i_output_module1[1:0]]), .Q(and10resu1_output_module1) );    

    MUX21X1 U3864(.IN1(ext_req_v_o[73:37][3]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+3]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][3]));
    MUX21X1 U3865(.IN1(ext_req_v_o[73:37][4]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+4]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][4]));
    MUX21X1 U3866(.IN1(ext_req_v_o[73:37][5]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+5]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][5]));
    MUX21X1 U3867(.IN1(ext_req_v_o[73:37][6]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+6]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][6]));
    MUX21X1 U3868(.IN1(ext_req_v_o[73:37][7]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+7]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][7]));
    MUX21X1 U3869(.IN1(ext_req_v_o[73:37][8]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+8]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][8]));
    MUX21X1 U3870(.IN1(ext_req_v_o[73:37][9]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+9]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][9]));
    MUX21X1 U3871(.IN1(ext_req_v_o[73:37][10]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+10]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][10]));
    MUX21X1 U3872(.IN1(ext_req_v_o[73:37][11]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+11]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][11]));
    MUX21X1 U3873(.IN1(ext_req_v_o[73:37][12]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+12]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][12]));
    MUX21X1 U3874(.IN1(ext_req_v_o[73:37][13]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+13]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][13]));
    MUX21X1 U3875(.IN1(ext_req_v_o[73:37][14]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+14]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][14]));
    MUX21X1 U3876(.IN1(ext_req_v_o[73:37][15]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+15]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][15]));
    MUX21X1 U3877(.IN1(ext_req_v_o[73:37][16]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+16]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][16]));
    MUX21X1 U3878(.IN1(ext_req_v_o[73:37][17]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+17]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][17]));
    MUX21X1 U3879(.IN1(ext_req_v_o[73:37][18]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+18]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][18]));
    MUX21X1 U3880(.IN1(ext_req_v_o[73:37][19]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+19]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][19]));
    MUX21X1 U3881(.IN1(ext_req_v_o[73:37][20]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+20]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][20]));
    MUX21X1 U3882(.IN1(ext_req_v_o[73:37][21]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+21]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][21]));
    MUX21X1 U3883(.IN1(ext_req_v_o[73:37][22]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+22]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][22]));
    MUX21X1 U3884(.IN1(ext_req_v_o[73:37][23]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+23]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][23]));
    MUX21X1 U3885(.IN1(ext_req_v_o[73:37][24]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+24]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][24]));
    MUX21X1 U3886(.IN1(ext_req_v_o[73:37][25]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+25]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][25]));
    MUX21X1 U3887(.IN1(ext_req_v_o[73:37][26]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+26]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][26]));
    MUX21X1 U3888(.IN1(ext_req_v_o[73:37][27]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+27]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][27]));
    MUX21X1 U3889(.IN1(ext_req_v_o[73:37][28]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+28]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][28]));
    MUX21X1 U3890(.IN1(ext_req_v_o[73:37][29]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+29]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][29]));
    MUX21X1 U3891(.IN1(ext_req_v_o[73:37][30]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+30]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][30]));
    MUX21X1 U3892(.IN1(ext_req_v_o[73:37][31]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+31]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][31]));
    MUX21X1 U3893(.IN1(ext_req_v_o[73:37][32]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+32]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][32]));
    MUX21X1 U3894(.IN1(ext_req_v_o[73:37][33]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+33]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][33]));
    MUX21X1 U3895(.IN1(ext_req_v_o[73:37][34]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+34]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][34]));
    MUX21X1 U3896(.IN1(ext_req_v_o[73:37][35]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+35]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][35]));
    MUX21X1 U3897(.IN1(ext_req_v_o[73:37][36]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37+36]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][36]));

    MUX21X1 U3898(.IN1(ext_req_v_o[73:37][0]), .IN2(int_map_req_v[184:148][i_output_module1[1:0]*37]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][0]);
    MUX21X1 U3899(.IN1(ext_req_v_o[73:37][1]), .IN2(vc_ch_act_out_output_module1[0]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][1]);
    MUX21X1 U3900(.IN1(ext_req_v_o[73:37][2]), .IN2(vc_ch_act_out_output_module1[1]), .S(and10resu1_output_module1) ,.Q(ext_req_v_o[73:37][2]);    
    MUX21X1 U3901(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3902(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b1), .S(and10resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    

    AND2X1 U3903 ( .IN1(and9resu1_output_module1), .IN2(nand1resu_output_module1), .Q(and11resu1_output_module1) );    
    MUX21X1 U3904(.IN1(_sv2v_jump_output_module1[0]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[0]);
    MUX21X1 U3905(.IN1(_sv2v_jump_output_module1[1]), .IN2(1'b0), .S(and11resu1_output_module1) ,.Q(_sv2v_jump_output_module1[1]);    
    
 





    BUFX1 U3906 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[0]) );
    BUFX1 U3907 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter122[1]) );
    BUFX1 U3908 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3909 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3910 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    XNOR2X1 U3911 ( .IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter122) );
    MUX21X1 U3912 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U3913 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    INVX1 U3914 ( .A(i_high_prior_arbiter122[0]), .Y(i_0_not_high_prior_arbiter122) );
    MUX21X1 U3915 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter122), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[0]);
    MUX21X1 U3916 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter122[0]), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(raw_grant[1]);
    MUX21X1 U3917 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U3918 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b1), .S(valid_from_im_output_module2[3:0][i_high_prior_arbiter122[0]]), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    NAND2X1 U3919 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(_sv2v_jump_high_prior_arbiter122[1]), .QN(nandres_high_prior_arbiter122) );
    MUX21X1 U3920 (.IN1(_sv2v_jump_high_prior_arbiter122[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[0]));
    MUX21X1 U3921 (.IN1(_sv2v_jump_high_prior_arbiter122[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter122), .Q(_sv2v_jump_high_prior_arbiter122[1]));
    HADDX1 U3922 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U3923 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );
    HADDX1 U3924 ( .A0(i_high_prior_arbiter122[0]), .B0(1'b1), .C1(i_high_prior_arbiter122[1]), .SO(i_high_prior_arbiter122[0]) );



    BUFX1 U3925 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[0]) );
    BUFX1 U3926 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter222[1]) );
    BUFX1 U3927 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3928 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3929 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    XNOR2X1 U3930 ( .IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter222) );
    MUX21X1 U3931 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U3932 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    INVX1 U3933 ( .A(i_high_prior_arbiter222[0]), .Y(i_0_not_high_prior_arbiter222) );
    MUX21X1 U3934 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter222), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[0]);
    MUX21X1 U3935 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter222[0]), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(masked_grant[1]);
    MUX21X1 U3936 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U3937 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter222[0]]), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    NAND2X1 U3938 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(_sv2v_jump_high_prior_arbiter222[1]), .QN(nandres_high_prior_arbiter222) );
    MUX21X1 U3939 (.IN1(_sv2v_jump_high_prior_arbiter222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[0]));
    MUX21X1 U3940 (.IN1(_sv2v_jump_high_prior_arbiter222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter222), .Q(_sv2v_jump_high_prior_arbiter222[1]));
    HADDX1 U3941 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U3942 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    HADDX1 U3943 ( .A0(i_high_prior_arbiter222[0]), .B0(1'b1), .C1(i_high_prior_arbiter222[1]), .SO(i_high_prior_arbiter222[0]) );
    

    BUFX1 U3944 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[0]) );
    BUFX1 U3945 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter22[1]) );
    AND2X1 U3946 ( .A(mask_ff_rr_arbiter22[0]), .B(valid_from_im_output_module2[3:0][0]), .Y(mask_req_rr_arbiter22[0]) );
    AND2X1 U3947 ( .A(mask_ff_rr_arbiter22[1]), .B(valid_from_im_output_module2[3:0][1]), .Y(mask_req_rr_arbiter22[1]) );
    BUFX1 U3948 ( .A(mask_ff_rr_arbiter22[0]), .Y(next_mask_rr_arbiter22[0]) );
    BUFX1 U3949 ( .A(mask_ff_rr_arbiter22[1]), .Y(next_mask_rr_arbiter22[1]) );
    XNOR2X1 U3950 ( .IN1(mask_req_rr_arbiter22[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter22) );
    XNOR2X1 U3951 ( .IN1(mask_req_rr_arbiter22[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter22) );
    MUX21X1 U3952 (.IN1(masked_grant_rr_arbiter22[0]), .IN2(raw_grant_rr_arbiter22[0]), .S(xnor0res_rr_arbiter22), .Q(grant_im_output_module2[3:0][0]));
    MUX21X1 U3953 (.IN1(masked_grant_rr_arbiter22[1]), .IN2(raw_grant_rr_arbiter22[1]), .S(xnor1res_rr_arbiter22), .Q(grant_im_output_module2[3:0][1]));

    BUFX1 U3954 ( .A(1'b0), .Y(i_rr_arbiter22[1]) );
    MUX21X1 U3955 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter22[0]));

    AND2X1 U3956 ( .A(_sv2v_jump_rr_rr_arbiter22[1]), .B(1'b0), .Y(firstif_rr_arbiter22) );
    MUX21X1 U3957 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U3958 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(firstif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    AND2X1 U3959 ( .A(firstif_rr_arbiter22), .B(grant_im_output_module2[3:0][i_rr_arbiter22[0]]), .Y(secondif_rr_arbiter22) );
    MUX21X1 U3960 (.IN1(next_mask_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[0]));
    MUX21X1 U3961 (.IN1(next_mask_rr_arbiter22[1]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(next_mask_rr_arbiter22[1]));
    MUX21X1 U3962 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter22[0]), .Q(j_rr_arbiter22[0]));
    AND2X1 U3963 ( .A(secondif_rr_arbiter22), .B(j_rr_arbiter22[0]), .Y(thirdif_rr_arbiter22) );
    MUX21X1 U3964 (.IN1(next_mask_rr_arbiter22[j_rr_arbiter22[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter22), .Q(next_mask_rr_arbiter22[j_rr_arbiter22[0]]));
    MUX21X1 U3965 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U3966 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b1), .S(secondif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));
    NAND2X1 U3967 ( .IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(_sv2v_jump_rr_rr_arbiter22[1]), .QN(fourthif_rr_arbiter22) );
    MUX21X1 U3968 (.IN1(_sv2v_jump_rr_rr_arbiter22[0]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[0]));
    MUX21X1 U3969 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(fourthif_rr_arbiter22), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    MUX21X1 U3970 (.IN1(_sv2v_jump_rr_rr_arbiter22[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter22[1]));

    DFFX2 U3971 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter22) );
    DFFX2 U3972 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter22) );
    MUX21X1 U3973 (.IN1(mask_ff_rr_arbiter22[0]), .IN2(next_mask_rr_arbiter22[0]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[0]));
    MUX21X1 U3974 (.IN1(mask_ff_rr_arbiter22[1]), .IN2(next_mask_rr_arbiter22[1]), .S(tail_flit_im_output_module2[0]), .Q(temp_mask_ff_rr_arbiter2222[1]));
    MUX21X1 U3975 (.IN1(temp_mask_ff_rr_arbiter2222), .IN2(1'sb1), .S(arst_value_rr_arbiter22), .Q(mask_ff_rr_arbiter22[0]));



    BUFX1 U3976 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[0]) );
    BUFX1 U3977 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1221[1]) );
    BUFX1 U3978 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U3979 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U3980 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    XNOR2X1 U3981 ( .IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1221) );
    MUX21X1 U3982 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U3983 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    INVX1 U3984 ( .A(i_high_prior_arbiter1221[0]), .Y(i_0_not_high_prior_arbiter1221) );
    MUX21X1 U3985 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1221), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[0]);
    MUX21X1 U3986 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1221[0]), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(raw_grant[1]);
    MUX21X1 U3987 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U3988 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b1), .S(valid_from_im_output_module2[7:4][i_high_prior_arbiter1221[0]]), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    NAND2X1 U3989 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(_sv2v_jump_high_prior_arbiter1221[1]), .QN(nandres_high_prior_arbiter1221) );
    MUX21X1 U3990 (.IN1(_sv2v_jump_high_prior_arbiter1221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[0]));
    MUX21X1 U3991 (.IN1(_sv2v_jump_high_prior_arbiter1221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1221), .Q(_sv2v_jump_high_prior_arbiter1221[1]));
    HADDX1 U3992 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U3993 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );
    HADDX1 U3994 ( .A0(i_high_prior_arbiter1221[0]), .B0(1'b1), .C1(i_high_prior_arbiter1221[1]), .SO(i_high_prior_arbiter1221[0]) );



    BUFX1 U3995 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[0]) );
    BUFX1 U3996 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2221[1]) );
    BUFX1 U3997 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U3998 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U3999 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    XNOR2X1 U4000 ( .IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter22212) );
    MUX21X1 U4001 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U4002 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    INVX1 U4003 ( .A(i_high_prior_arbiter2221[0]), .Y(i_0_not_high_prior_arbiter22212) );
    MUX21X1 U4004 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter22212), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[0]);
    MUX21X1 U4005 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2221[0]), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(masked_grant[1]);
    MUX21X1 U4006 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U4007 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2221[0]]), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    NAND2X1 U4008 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(_sv2v_jump_high_prior_arbiter2221[1]), .QN(nandres_high_prior_arbiter22212) );
    MUX21X1 U4009 (.IN1(_sv2v_jump_high_prior_arbiter2221[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[0]));
    MUX21X1 U4010 (.IN1(_sv2v_jump_high_prior_arbiter2221[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter22212), .Q(_sv2v_jump_high_prior_arbiter2221[1]));
    HADDX1 U4011 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U4012 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    HADDX1 U4013 ( .A0(i_high_prior_arbiter2221[0]), .B0(1'b1), .C1(i_high_prior_arbiter2221[1]), .SO(i_high_prior_arbiter2221[0]) );
    

    BUFX1 U4014 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[0]) );
    BUFX1 U4015 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter221[1]) );
    AND2X1 U4016 ( .A(mask_ff_rr_arbiter221[0]), .B(valid_from_im_output_module2[7:4][0]), .Y(mask_req_rr_arbiter221[0]) );
    AND2X1 U4017 ( .A(mask_ff_rr_arbiter221[1]), .B(valid_from_im_output_module2[7:4][1]), .Y(mask_req_rr_arbiter221[1]) );
    BUFX1 U4018 ( .A(mask_ff_rr_arbiter221[0]), .Y(next_mask_rr_arbiter221[0]) );
    BUFX1 U4019 ( .A(mask_ff_rr_arbiter221[1]), .Y(next_mask_rr_arbiter221[1]) );
    XNOR2X1 U4020 ( .IN1(mask_req_rr_arbiter221[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter221) );
    XNOR2X1 U4021 ( .IN1(mask_req_rr_arbiter221[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter221) );
    MUX21X1 U4022 (.IN1(masked_grant_rr_arbiter221[0]), .IN2(raw_grant_rr_arbiter221[0]), .S(xnor0res_rr_arbiter221), .Q(grant_im_output_module2[7:4][0]));
    MUX21X1 U4023 (.IN1(masked_grant_rr_arbiter221[1]), .IN2(raw_grant_rr_arbiter221[1]), .S(xnor1res_rr_arbiter221), .Q(grant_im_output_module2[7:4][1]));

    BUFX1 U4024 ( .A(1'b0), .Y(i_rr_arbiter221[1]) );
    MUX21X1 U4025 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter221[0]));

    AND2X1 U4026 ( .A(_sv2v_jump_rr_rr_arbiter221[1]), .B(1'b0), .Y(firstif_rr_arbiter221) );
    MUX21X1 U4027 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U4028 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(firstif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    AND2X1 U4029 ( .A(firstif_rr_arbiter221), .B(grant_im_output_module2[7:4][i_rr_arbiter221[0]]), .Y(secondif_rr_arbiter221) );
    MUX21X1 U4030 (.IN1(next_mask_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[0]));
    MUX21X1 U4031 (.IN1(next_mask_rr_arbiter221[1]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(next_mask_rr_arbiter221[1]));
    MUX21X1 U4032 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter221[0]), .Q(j_rr_arbiter221[0]));
    AND2X1 U4033 ( .A(secondif_rr_arbiter221), .B(j_rr_arbiter221[0]), .Y(thirdif_rr_arbiter221) );
    MUX21X1 U4034 (.IN1(next_mask_rr_arbiter221[j_rr_arbiter221[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter221), .Q(next_mask_rr_arbiter221[j_rr_arbiter221[0]]));
    MUX21X1 U4035 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U4036 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b1), .S(secondif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));
    NAND2X1 U4037 ( .IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(_sv2v_jump_rr_rr_arbiter221[1]), .QN(fourthif_rr_arbiter221) );
    MUX21X1 U4038 (.IN1(_sv2v_jump_rr_rr_arbiter221[0]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[0]));
    MUX21X1 U4039 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(fourthif_rr_arbiter221), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    MUX21X1 U4040 (.IN1(_sv2v_jump_rr_rr_arbiter221[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter221[1]));

    DFFX2 U4041 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter221) );
    DFFX2 U4042 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter221) );
    MUX21X1 U4043 (.IN1(mask_ff_rr_arbiter221[0]), .IN2(next_mask_rr_arbiter221[0]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[0]));
    MUX21X1 U4044 (.IN1(mask_ff_rr_arbiter221[1]), .IN2(next_mask_rr_arbiter221[1]), .S(tail_flit_im_output_module2[1]), .Q(temp_mask_ff_rr_arbiter222211[1]));
    MUX21X1 U4045 (.IN1(temp_mask_ff_rr_arbiter222211), .IN2(1'sb1), .S(arst_value_rr_arbiter221), .Q(mask_ff_rr_arbiter221[0]));





    BUFX1 U4046 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[0]) );
    BUFX1 U4047 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter1222[1]) );
    BUFX1 U4048 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4049 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4050 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    XNOR2X1 U4051 ( .IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter1222) );
    MUX21X1 U4052 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U4053 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    INVX1 U4054 ( .A(i_high_prior_arbiter1222[0]), .Y(i_0_not_high_prior_arbiter1222) );
    MUX21X1 U4055 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter1222), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[0]);
    MUX21X1 U4056 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter1222[0]), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(raw_grant[1]);
    MUX21X1 U4057 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U4058 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b1), .S(valid_from_im_output_module2[11:8][i_high_prior_arbiter1222[0]]), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    NAND2X1 U4059 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(_sv2v_jump_high_prior_arbiter1222[1]), .QN(nandres_high_prior_arbiter1222) );
    MUX21X1 U4060 (.IN1(_sv2v_jump_high_prior_arbiter1222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[0]));
    MUX21X1 U4061 (.IN1(_sv2v_jump_high_prior_arbiter1222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter1222), .Q(_sv2v_jump_high_prior_arbiter1222[1]));
    HADDX1 U4062 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U4063 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );
    HADDX1 U4064 ( .A0(i_high_prior_arbiter1222[0]), .B0(1'b1), .C1(i_high_prior_arbiter1222[1]), .SO(i_high_prior_arbiter1222[0]) );



    BUFX1 U4065 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[0]) );
    BUFX1 U4066 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter2222[1]) );
    BUFX1 U4067 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4068 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4069 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    XNOR2X1 U4070 ( .IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2222) );
    MUX21X1 U4071 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U4072 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    INVX1 U4073 ( .A(i_high_prior_arbiter2222[0]), .Y(i_0_not_high_prior_arbiter2222) );
    MUX21X1 U4074 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2222), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[0]);
    MUX21X1 U4075 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter2222[0]), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(masked_grant[1]);
    MUX21X1 U4076 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U4077 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter2222[0]]), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    NAND2X1 U4078 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(_sv2v_jump_high_prior_arbiter2222[1]), .QN(nandres_high_prior_arbiter2222) );
    MUX21X1 U4079 (.IN1(_sv2v_jump_high_prior_arbiter2222[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[0]));
    MUX21X1 U4080 (.IN1(_sv2v_jump_high_prior_arbiter2222[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2222), .Q(_sv2v_jump_high_prior_arbiter2222[1]));
    HADDX1 U4081 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U4082 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    HADDX1 U4083 ( .A0(i_high_prior_arbiter2222[0]), .B0(1'b1), .C1(i_high_prior_arbiter2222[1]), .SO(i_high_prior_arbiter2222[0]) );
    

    BUFX1 U4084 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[0]) );
    BUFX1 U4085 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter222[1]) );
    AND2X1 U4086 ( .A(mask_ff_rr_arbiter222[0]), .B(valid_from_im_output_module2[11:8][0]), .Y(mask_req_rr_arbiter222[0]) );
    AND2X1 U4087 ( .A(mask_ff_rr_arbiter222[1]), .B(valid_from_im_output_module2[11:8][1]), .Y(mask_req_rr_arbiter222[1]) );
    BUFX1 U4088 ( .A(mask_ff_rr_arbiter222[0]), .Y(next_mask_rr_arbiter222[0]) );
    BUFX1 U4089 ( .A(mask_ff_rr_arbiter222[1]), .Y(next_mask_rr_arbiter222[1]) );
    XNOR2X1 U4090 ( .IN1(mask_req_rr_arbiter222[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter222) );
    XNOR2X1 U4091 ( .IN1(mask_req_rr_arbiter222[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter222) );
    MUX21X1 U4092 (.IN1(masked_grant_rr_arbiter222[0]), .IN2(raw_grant_rr_arbiter222[0]), .S(xnor0res_rr_arbiter222), .Q(grant_im_output_module2[11:8][0]));
    MUX21X1 U4093 (.IN1(masked_grant_rr_arbiter222[1]), .IN2(raw_grant_rr_arbiter222[1]), .S(xnor1res_rr_arbiter222), .Q(grant_im_output_module2[11:8][1]));

    BUFX1 U4094 ( .A(1'b0), .Y(i_rr_arbiter222[1]) );
    MUX21X1 U4095 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter222[0]));

    AND2X1 U4096 ( .A(_sv2v_jump_rr_rr_arbiter222[1]), .B(1'b0), .Y(firstif_rr_arbiter222) );
    MUX21X1 U4097 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U4098 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(firstif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    AND2X1 U4099 ( .A(firstif_rr_arbiter222), .B(grant_im_output_module2[11:8][i_rr_arbiter222[0]]), .Y(secondif_rr_arbiter222) );
    MUX21X1 U4100 (.IN1(next_mask_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[0]));
    MUX21X1 U4101 (.IN1(next_mask_rr_arbiter222[1]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(next_mask_rr_arbiter222[1]));
    MUX21X1 U4102 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter222[0]), .Q(j_rr_arbiter222[0]));
    AND2X1 U4103 ( .A(secondif_rr_arbiter222), .B(j_rr_arbiter222[0]), .Y(thirdif_rr_arbiter222) );
    MUX21X1 U4104 (.IN1(next_mask_rr_arbiter222[j_rr_arbiter222[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter222), .Q(next_mask_rr_arbiter222[j_rr_arbiter222[0]]));
    MUX21X1 U4105 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U4106 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b1), .S(secondif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));
    NAND2X1 U4107 ( .IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(_sv2v_jump_rr_rr_arbiter222[1]), .QN(fourthif_rr_arbiter222) );
    MUX21X1 U4108 (.IN1(_sv2v_jump_rr_rr_arbiter222[0]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[0]));
    MUX21X1 U4109 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(fourthif_rr_arbiter222), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    MUX21X1 U4110 (.IN1(_sv2v_jump_rr_rr_arbiter222[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter222[1]));

    DFFX2 U4111 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter222) );
    DFFX2 U4112 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter222) );
    MUX21X1 U4113 (.IN1(mask_ff_rr_arbiter222[0]), .IN2(next_mask_rr_arbiter222[0]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[0]));
    MUX21X1 U4114 (.IN1(mask_ff_rr_arbiter222[1]), .IN2(next_mask_rr_arbiter222[1]), .S(tail_flit_im_output_module2[2]), .Q(temp_mask_ff_rr_arbiter222222[1]));
    MUX21X1 U4115 (.IN1(temp_mask_ff_rr_arbiter222222), .IN2(1'sb1), .S(arst_value_rr_arbiter222), .Q(mask_ff_rr_arbiter222[0]));


    XNOR2X1 U4116 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37]), .IN2(vc_channel_output_module2[1]), .QN(xnor1resu1_output_module2) );
    XNOR2X1 U4117 ( .IN1(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37-1]), .IN2(vc_channel_output_module2[0]), .QN(xnor2resu1_output_module2) );
    AND2X1 U4118 ( .IN1(xnor1resu1_output_module2), .IN2(xnor2resu1_output_module2), .Q(and1resu1_output_module2) );
    MUX21X1 U4119 (.IN1(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]), .IN2(1'b1), .S(and1resu1_output_module2), .Q(valid_from_im_output_module2[(vc_channel_output_module2[1:0]*4) + in_mod_output_module2[1:0]]);
    HADDX1 U4120 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4121 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4122 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4123 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4124 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4125 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4126 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4127 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4128 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4129 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );  
    HADDX1 U4130 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4131 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4132 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4133 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) ); 
    XOR2X1 U4134 ( .IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .Q(xor1resu1_output_module2) );
    MUX21X1 U4135 (.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[0]));
    MUX21X1 U4136 (.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2[1]));
    MUX21X1 U4137 (.IN1(_sv2v_jump_output_module2_1[0]), .IN2(_sv2v_jump_output_module2[0]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[0]));
    MUX21X1 U4138 (.IN1(_sv2v_jump_output_module2_1[1]), .IN2(_sv2v_jump_output_module2[1]), .S(xor1resu1_output_module2), .Q(_sv2v_jump_output_module2_1[1]));
    AND2X1 U4139 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[vc_channel_output_module2[1:0]*4+in_mod_output_module2[1:0]]), .Q(and2resu1_output_module2) );

    MUX21X1 U4140(.IN1(head_flit_output_module2[3]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+3]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[3]));
    MUX21X1 U4141(.IN1(head_flit_output_module2[4]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+4]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[4]));
    MUX21X1 U4142(.IN1(head_flit_output_module2[5]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+5]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[5]));
    MUX21X1 U4143(.IN1(head_flit_output_module2[6]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+6]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[6]));
    MUX21X1 U4144(.IN1(head_flit_output_module2[7]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+7]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[7]));
    MUX21X1 U4145(.IN1(head_flit_output_module2[8]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+8]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[8]));
    MUX21X1 U4146(.IN1(head_flit_output_module2[9]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+9]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[9]));
    MUX21X1 U4147(.IN1(head_flit_output_module2[10]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+10]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[10]));
    MUX21X1 U4148(.IN1(head_flit_output_module2[11]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+11]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[11]));
    MUX21X1 U4149(.IN1(head_flit_output_module2[12]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+12]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[12]));
    MUX21X1 U4150(.IN1(head_flit_output_module2[13]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+13]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[13]));
    MUX21X1 U4151(.IN1(head_flit_output_module2[14]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+14]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[14]));
    MUX21X1 U4152(.IN1(head_flit_output_module2[15]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+15]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[15]));
    MUX21X1 U4153(.IN1(head_flit_output_module2[16]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+16]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[16]));
    MUX21X1 U4154(.IN1(head_flit_output_module2[17]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+17]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[17]));
    MUX21X1 U4155(.IN1(head_flit_output_module2[18]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+18]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[18]));
    MUX21X1 U4156(.IN1(head_flit_output_module2[19]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+19]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[19]));
    MUX21X1 U4157(.IN1(head_flit_output_module2[20]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+20]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[20]));
    MUX21X1 U4158(.IN1(head_flit_output_module2[21]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+21]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[21]));
    MUX21X1 U4159(.IN1(head_flit_output_module2[22]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+22]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[22]));
    MUX21X1 U4160(.IN1(head_flit_output_module2[23]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+23]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[23]));
    MUX21X1 U4161(.IN1(head_flit_output_module2[24]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+24]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[24]));
    MUX21X1 U4162(.IN1(head_flit_output_module2[25]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+25]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[25]));
    MUX21X1 U4163(.IN1(head_flit_output_module2[26]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+26]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[26]));
    MUX21X1 U4164(.IN1(head_flit_output_module2[27]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+27]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[27]));
    MUX21X1 U4165(.IN1(head_flit_output_module2[28]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+28]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[28]));
    MUX21X1 U4166(.IN1(head_flit_output_module2[29]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+29]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[29]));
    MUX21X1 U4167(.IN1(head_flit_output_module2[30]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+30]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[30]));
    MUX21X1 U4168(.IN1(head_flit_output_module2[31]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+31]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[31]));
    MUX21X1 U4169(.IN1(head_flit_output_module2[32]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+32]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[32]));
    MUX21X1 U4170(.IN1(head_flit_output_module2[33]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+33]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[33]));
    MUX21X1 U4171(.IN1(head_flit_output_module2[34]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+34]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[34]));
    MUX21X1 U4172(.IN1(head_flit_output_module2[35]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+35]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[35]));
    MUX21X1 U4173(.IN1(head_flit_output_module2[36]), .IN2(nt_map_req_v[332:296][in_mod_output_module2[1:0]*37+36]), .S(and2resu1_output_module2) ,.Q(head_flit_output_module2[36]));

    INVX1 U4174 ( .A(head_flit_output_module2[32]), .Y(head_flit_output_module2_32_not_output_module2) );
    AND2X1 U4175 ( .IN1(head_flit_output_module2_32_not_output_module2), .IN2(head_flit_output_module2[33]), .Q(and3resu1_output_module2) );
    NOR4X1 U4176 (.IN1(head_flit_output_module2[29]), .IN2(head_flit_output_module2[28]), .IN3(head_flit_output_module2[27]), .IN4(head_flit_output_module2[26]), .Q(nor23resu1_output_module2) );
    NOR4X1 U4177 (.IN1(head_flit_output_module2[25]), .IN2(head_flit_output_module2[24]), .IN3(head_flit_output_module2[23]), .IN4(head_flit_output_module2[22]), .Q(nor23resu2_output_module2) );
    AND2X1 U4178 ( .IN1(nor23resu1_output_module2), .IN2(nor23resu2_output_module2), .Q(and4resu1_output_module2) );
    NOR2X1 U4179 (.IN1(head_flit_output_module2[33]), .IN2(head_flit_output_module2[32]), .Q(nor23resu3_output_module2) );
    AND2X1 U4180 ( .IN1(nor23resu3_output_module2), .IN2(and4resu1_output_module2), .Q(and5resu1_output_module2) );    
    OR2X1 U4181 (.IN1(and3resu1_output_module2), .IN2(nor23resu3_output_module2), .Q(or12resu12_output_module2) );
    AND2X1 U4182 ( .IN1(ext_resp_v_i[3:2][0]), .IN2(or12resu12_output_module2), .Q(and6resu1_output_module2) );    
    MUX21X1 U4183(.IN1(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]), .IN2(and6resu1_output_module2), .S(and2resu1_output_module2) ,.Q(tail_flit_im_output_module2[vc_channel_output_module2[1:0]]);
    MUX21X1 U4184(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4185(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and2resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    NAND2X1 U4186(.A(_sv2v_jump_output_module2[0]),.B(_sv2v_jump_output_module2[1]),.Y(nand1resu_output_module2));

    AND2X1 U4187 ( .IN1(xor1resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and7resu1) );    
    MUX21X1 U4188(.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4189(.IN1(_sv2v_jump_output_module2[1]), .IN2(_sv2v_jump_output_module2_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    MUX21X1 U4190(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4191(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module2[1]);

    HADDX1 U4192 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4193 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4194 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4195 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4196 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4197 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4198 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4199 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4200 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4201 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4202 ( .A0(vc_channel_output_module2[0]), .B0(1'b1), .C1(vc_channel_output_module2[1]), .SO(vc_channel_output_module2[0]) );
    HADDX1 U4203 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4204 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4205 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );
    HADDX1 U4206 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(in_mod_output_module2[1]), .SO(in_mod_output_module2[0]) );



    BUFX1 U4207(.A(1'b0), .Y(_sv2v_jump_output_module2[0]));
    BUFX1 U4208(.A(1'b0), .Y(_sv2v_jump_output_module2[1]));
    AND2X1 U4209 ( .IN1(xor1resu1_output_module2), .IN2(grant_im_output_module2[i_output_module2[1:0] * 4+:4]), .Q(and8resu1_output_module2) );    
    MUX21X1 U4210(.IN1(vc_ch_act_out_output_module2[0]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[0]);
    MUX21X1 U4211(.IN1(vc_ch_act_out_output_module2[1]), .IN2(i_output_module2[1:0]), .S(and8resu1_output_module2) ,.Q(vc_ch_act_out_output_module2[1]);
    MUX21X1 U4212(.IN1(req_out_output_module2), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(req_out_output_module2);
    MUX21X1 U4213(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4214(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and8resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);
    HADDX1 U4215 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U4216 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    HADDX1 U4217 ( .A0(in_mod_output_module2[0]), .B0(1'b1), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );

    NOR2X1 U4218 (.IN1(_sv2v_jump_output_module2[0]), .IN2(_sv2v_jump_output_module2[1]), .Q(norfinresu1_output_module2) );
    AND2X1 U4219 ( .IN1(norfinresu1_output_module2), .IN2(req_out_output_module2), .Q(and9resu1_output_module2) );    
    HADDX1 U4220 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module2[1]), .SO(i_output_module2[0]) );
    AND2X1 U4221 ( .IN1(and9resu1_output_module2), .IN2(grant_im_output_module2[(vc_ch_act_out_output_module2 * 4) + i_output_module2[1:0]]), .Q(and10resu1_output_module2) );    

    MUX21X1 U4222(.IN1(ext_req_v_o[110:74][3]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+3]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][3]));
    MUX21X1 U4223(.IN1(ext_req_v_o[110:74][4]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+4]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][4]));
    MUX21X1 U4224(.IN1(ext_req_v_o[110:74][5]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+5]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][5]));
    MUX21X1 U4225(.IN1(ext_req_v_o[110:74][6]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+6]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][6]));
    MUX21X1 U4226(.IN1(ext_req_v_o[110:74][7]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+7]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][7]));
    MUX21X1 U4227(.IN1(ext_req_v_o[110:74][8]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+8]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][8]));
    MUX21X1 U4228(.IN1(ext_req_v_o[110:74][9]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+9]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][9]));
    MUX21X1 U4229(.IN1(ext_req_v_o[110:74][10]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+10]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][10]));
    MUX21X1 U4230(.IN1(ext_req_v_o[110:74][11]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+11]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][11]));
    MUX21X1 U4231(.IN1(ext_req_v_o[110:74][12]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+12]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][12]));
    MUX21X1 U4232(.IN1(ext_req_v_o[110:74][13]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+13]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][13]));
    MUX21X1 U4233(.IN1(ext_req_v_o[110:74][14]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+14]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][14]));
    MUX21X1 U4234(.IN1(ext_req_v_o[110:74][15]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+15]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][15]));
    MUX21X1 U4235(.IN1(ext_req_v_o[110:74][16]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+16]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][16]));
    MUX21X1 U4236(.IN1(ext_req_v_o[110:74][17]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+17]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][17]));
    MUX21X1 U4237(.IN1(ext_req_v_o[110:74][18]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+18]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][18]));
    MUX21X1 U4238(.IN1(ext_req_v_o[110:74][19]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+19]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][19]));
    MUX21X1 U4239(.IN1(ext_req_v_o[110:74][20]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+20]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][20]));
    MUX21X1 U4240(.IN1(ext_req_v_o[110:74][21]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+21]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][21]));
    MUX21X1 U4241(.IN1(ext_req_v_o[110:74][22]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+22]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][22]));
    MUX21X1 U4242(.IN1(ext_req_v_o[110:74][23]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+23]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][23]));
    MUX21X1 U4243(.IN1(ext_req_v_o[110:74][24]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+24]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][24]));
    MUX21X1 U4244(.IN1(ext_req_v_o[110:74][25]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+25]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][25]));
    MUX21X1 U4245(.IN1(ext_req_v_o[110:74][26]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+26]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][26]));
    MUX21X1 U4246(.IN1(ext_req_v_o[110:74][27]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+27]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][27]));
    MUX21X1 U4247(.IN1(ext_req_v_o[110:74][28]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+28]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][28]));
    MUX21X1 U4248(.IN1(ext_req_v_o[110:74][29]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+29]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][29]));
    MUX21X1 U4249(.IN1(ext_req_v_o[110:74][30]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+30]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][30]));
    MUX21X1 U4250(.IN1(ext_req_v_o[110:74][31]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+31]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][31]));
    MUX21X1 U4251(.IN1(ext_req_v_o[110:74][32]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+32]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][32]));
    MUX21X1 U4252(.IN1(ext_req_v_o[110:74][33]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+33]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][33]));
    MUX21X1 U4253(.IN1(ext_req_v_o[110:74][34]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+34]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][34]));
    MUX21X1 U4254(.IN1(ext_req_v_o[110:74][35]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+35]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][35]));
    MUX21X1 U4255(.IN1(ext_req_v_o[110:74][36]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37+36]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][36]));

    MUX21X1 U4256(.IN1(ext_req_v_o[110:74][0]), .IN2(nt_map_req_v[332:296][i_output_module2[1:0]*37]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][0]);
    MUX21X1 U4257(.IN1(ext_req_v_o[110:74][1]), .IN2(vc_ch_act_out_output_module2[0]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][1]);
    MUX21X1 U4258(.IN1(ext_req_v_o[110:74][2]), .IN2(vc_ch_act_out_output_module2[1]), .S(and10resu1_output_module2) ,.Q(ext_req_v_o[110:74][2]);    
    MUX21X1 U4259(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4260(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b1), .S(and10resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);    

    AND2X1 U4261 ( .IN1(and9resu1_output_module2), .IN2(nand1resu_output_module2), .Q(and11resu1_output_module2) );    
    MUX21X1 U4262(.IN1(_sv2v_jump_output_module2[0]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[0]);
    MUX21X1 U4263(.IN1(_sv2v_jump_output_module2[1]), .IN2(1'b0), .S(and11resu1_output_module2) ,.Q(_sv2v_jump_output_module2[1]);   










    BUFX1 U4264 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[0]) );
    BUFX1 U4265 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter13[1]) );
    BUFX1 U4266 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4267 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4268 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    XNOR2X1 U4269 ( .IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter13) );
    MUX21X1 U4270 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U4271 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    INVX1 U4272 ( .A(i_high_prior_arbiter13[0]), .Y(i_0_not_high_prior_arbiter13) );
    MUX21X1 U4273 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter13), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[0]);
    MUX21X1 U4274 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter13[0]), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(raw_grant[1]);
    MUX21X1 U4275 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U4276 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b1), .S(valid_from_im_output_module3[3:0][i_high_prior_arbiter13[0]]), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    NAND2X1 U4277 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(_sv2v_jump_high_prior_arbiter13[1]), .QN(nandres_high_prior_arbiter13) );
    MUX21X1 U4278 (.IN1(_sv2v_jump_high_prior_arbiter13[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[0]));
    MUX21X1 U4279 (.IN1(_sv2v_jump_high_prior_arbiter13[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter13), .Q(_sv2v_jump_high_prior_arbiter13[1]));
    HADDX1 U4280 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U4281 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );
    HADDX1 U4282 ( .A0(i_high_prior_arbiter13[0]), .B0(1'b1), .C1(i_high_prior_arbiter13[1]), .SO(i_high_prior_arbiter13[0]) );



    BUFX1 U4283 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[0]) );
    BUFX1 U4284 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter23[1]) );
    BUFX1 U4285 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4286 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4287 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    XNOR2X1 U4288 ( .IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter23) );
    MUX21X1 U4289 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U4290 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    INVX1 U4291 ( .A(i_high_prior_arbiter23[0]), .Y(i_0_not_high_prior_arbiter23) );
    MUX21X1 U4292 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter23), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[0]);
    MUX21X1 U4293 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter23[0]), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(masked_grant[1]);
    MUX21X1 U4294 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U4295 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter23[0]]), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    NAND2X1 U4296 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(_sv2v_jump_high_prior_arbiter23[1]), .QN(nandres_high_prior_arbiter23) );
    MUX21X1 U4297 (.IN1(_sv2v_jump_high_prior_arbiter23[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[0]));
    MUX21X1 U4298 (.IN1(_sv2v_jump_high_prior_arbiter23[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter23), .Q(_sv2v_jump_high_prior_arbiter23[1]));
    HADDX1 U4299 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U4300 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    HADDX1 U4301 ( .A0(i_high_prior_arbiter23[0]), .B0(1'b1), .C1(i_high_prior_arbiter23[1]), .SO(i_high_prior_arbiter23[0]) );
    

    BUFX1 U4302 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[0]) );
    BUFX1 U4303 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter3[1]) );
    AND2X1 U4304 ( .A(mask_ff_rr_arbiter3[0]), .B(valid_from_im_output_module3[3:0][0]), .Y(mask_req_rr_arbiter3[0]) );
    AND2X1 U4305 ( .A(mask_ff_rr_arbiter3[1]), .B(valid_from_im_output_module3[3:0][1]), .Y(mask_req_rr_arbiter3[1]) );
    BUFX1 U4306 ( .A(mask_ff_rr_arbiter3[0]), .Y(next_mask_rr_arbiter3[0]) );
    BUFX1 U4307 ( .A(mask_ff_rr_arbiter3[1]), .Y(next_mask_rr_arbiter3[1]) );
    XNOR2X1 U4308 ( .IN1(mask_req_rr_arbiter3[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter3) );
    XNOR2X1 U4309 ( .IN1(mask_req_rr_arbiter3[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter3) );
    MUX21X1 U4310 (.IN1(masked_grant_rr_arbiter3[0]), .IN2(raw_grant_rr_arbiter3[0]), .S(xnor0res_rr_arbiter3), .Q(grant_im_output_module3[3:0][0]));
    MUX21X1 U4311 (.IN1(masked_grant_rr_arbiter3[1]), .IN2(raw_grant_rr_arbiter3[1]), .S(xnor1res_rr_arbiter3), .Q(grant_im_output_module3[3:0][1]));

    BUFX1 U4312 ( .A(1'b0), .Y(i_rr_arbiter3[1]) );
    MUX21X1 U4313 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter3[0]));

    AND2X1 U4314 ( .A(_sv2v_jump_rr_rr_arbiter3[1]), .B(1'b0), .Y(firstif_rr_arbiter3) );
    MUX21X1 U4315 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U4316 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(firstif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    AND2X1 U4317 ( .A(firstif_rr_arbiter3), .B(grant_im_output_module3[3:0][i_rr_arbiter3[0]]), .Y(secondif_rr_arbiter3) );
    MUX21X1 U4318 (.IN1(next_mask_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[0]));
    MUX21X1 U4319 (.IN1(next_mask_rr_arbiter3[1]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(next_mask_rr_arbiter3[1]));
    MUX21X1 U4320 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter3[0]), .Q(j_rr_arbiter3[0]));
    AND2X1 U4321 ( .A(secondif_rr_arbiter3), .B(j_rr_arbiter3[0]), .Y(thirdif_rr_arbiter3) );
    MUX21X1 U4322 (.IN1(next_mask_rr_arbiter3[j_rr_arbiter3[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter3), .Q(next_mask_rr_arbiter3[j_rr_arbiter3[0]]));
    MUX21X1 U4323 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U4324 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b1), .S(secondif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));
    NAND2X1 U4325 ( .IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(_sv2v_jump_rr_rr_arbiter3[1]), .QN(fourthif_rr_arbiter3) );
    MUX21X1 U4326 (.IN1(_sv2v_jump_rr_rr_arbiter3[0]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[0]));
    MUX21X1 U4327 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(fourthif_rr_arbiter3), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    MUX21X1 U4328 (.IN1(_sv2v_jump_rr_rr_arbiter3[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter3[1]));

    DFFX2 U4329 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter3) );
    DFFX2 U4330 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter3) );
    MUX21X1 U4331 (.IN1(mask_ff_rr_arbiter3[0]), .IN2(next_mask_rr_arbiter3[0]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[0]));
    MUX21X1 U4332 (.IN1(mask_ff_rr_arbiter3[1]), .IN2(next_mask_rr_arbiter3[1]), .S(tail_flit_im_output_module3[0]), .Q(temp_mask_ff_rr_arbiter33[1]));
    MUX21X1 U4333 (.IN1(temp_mask_ff_rr_arbiter33), .IN2(1'sb1), .S(arst_value_rr_arbiter3), .Q(mask_ff_rr_arbiter3[0]));



    BUFX1 U4334 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[0]) );
    BUFX1 U4335 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter131[1]) );
    BUFX1 U4336 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4337 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4338 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    XNOR2X1 U4339 ( .IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter131) );
    MUX21X1 U4340 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U4341 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    INVX1 U4342 ( .A(i_high_prior_arbiter131[0]), .Y(i_0_not_high_prior_arbiter131) );
    MUX21X1 U4343 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter131), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[0]);
    MUX21X1 U4344 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter131[0]), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(raw_grant[1]);
    MUX21X1 U4345 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U4346 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b1), .S(valid_from_im_output_module3[7:4][i_high_prior_arbiter131[0]]), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    NAND2X1 U4347 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(_sv2v_jump_high_prior_arbiter131[1]), .QN(nandres_high_prior_arbiter131) );
    MUX21X1 U4348 (.IN1(_sv2v_jump_high_prior_arbiter131[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[0]));
    MUX21X1 U4349 (.IN1(_sv2v_jump_high_prior_arbiter131[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter131), .Q(_sv2v_jump_high_prior_arbiter131[1]));
    HADDX1 U4350 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U4351 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );
    HADDX1 U4352 ( .A0(i_high_prior_arbiter131[0]), .B0(1'b1), .C1(i_high_prior_arbiter131[1]), .SO(i_high_prior_arbiter131[0]) );



    BUFX1 U4353 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[0]) );
    BUFX1 U4354 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter231[1]) );
    BUFX1 U4355 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4356 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4357 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    XNOR2X1 U4358 ( .IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2313) );
    MUX21X1 U4359 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U4360 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    INVX1 U4361 ( .A(i_high_prior_arbiter231[0]), .Y(i_0_not_high_prior_arbiter2313) );
    MUX21X1 U4362 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2313), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[0]);
    MUX21X1 U4363 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter231[0]), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(masked_grant[1]);
    MUX21X1 U4364 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U4365 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter231[0]]), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    NAND2X1 U4366 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(_sv2v_jump_high_prior_arbiter231[1]), .QN(nandres_high_prior_arbiter2313) );
    MUX21X1 U4367 (.IN1(_sv2v_jump_high_prior_arbiter231[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[0]));
    MUX21X1 U4368 (.IN1(_sv2v_jump_high_prior_arbiter231[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2313), .Q(_sv2v_jump_high_prior_arbiter231[1]));
    HADDX1 U4369 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U4370 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    HADDX1 U4371 ( .A0(i_high_prior_arbiter231[0]), .B0(1'b1), .C1(i_high_prior_arbiter231[1]), .SO(i_high_prior_arbiter231[0]) );
    

    BUFX1 U4372 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[0]) );
    BUFX1 U4373 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter31[1]) );
    AND2X1 U4374 ( .A(mask_ff_rr_arbiter31[0]), .B(valid_from_im_output_module3[7:4][0]), .Y(mask_req_rr_arbiter31[0]) );
    AND2X1 U4375 ( .A(mask_ff_rr_arbiter31[1]), .B(valid_from_im_output_module3[7:4][1]), .Y(mask_req_rr_arbiter31[1]) );
    BUFX1 U4376 ( .A(mask_ff_rr_arbiter31[0]), .Y(next_mask_rr_arbiter31[0]) );
    BUFX1 U4377 ( .A(mask_ff_rr_arbiter31[1]), .Y(next_mask_rr_arbiter31[1]) );
    XNOR2X1 U4378 ( .IN1(mask_req_rr_arbiter31[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter31) );
    XNOR2X1 U4379 ( .IN1(mask_req_rr_arbiter31[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter31) );
    MUX21X1 U4380 (.IN1(masked_grant_rr_arbiter31[0]), .IN2(raw_grant_rr_arbiter31[0]), .S(xnor0res_rr_arbiter31), .Q(grant_im_output_module3[7:4][0]));
    MUX21X1 U4381 (.IN1(masked_grant_rr_arbiter31[1]), .IN2(raw_grant_rr_arbiter31[1]), .S(xnor1res_rr_arbiter31), .Q(grant_im_output_module3[7:4][1]));

    BUFX1 U4382 ( .A(1'b0), .Y(i_rr_arbiter31[1]) );
    MUX21X1 U4383 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter31[0]));

    AND2X1 U4384 ( .A(_sv2v_jump_rr_rr_arbiter31[1]), .B(1'b0), .Y(firstif_rr_arbiter31) );
    MUX21X1 U4385 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U4386 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(firstif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    AND2X1 U4387 ( .A(firstif_rr_arbiter31), .B(grant_im_output_module3[7:4][i_rr_arbiter31[0]]), .Y(secondif_rr_arbiter31) );
    MUX21X1 U4388 (.IN1(next_mask_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[0]));
    MUX21X1 U4389 (.IN1(next_mask_rr_arbiter31[1]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(next_mask_rr_arbiter31[1]));
    MUX21X1 U4390 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter31[0]), .Q(j_rr_arbiter31[0]));
    AND2X1 U4391 ( .A(secondif_rr_arbiter31), .B(j_rr_arbiter31[0]), .Y(thirdif_rr_arbiter31) );
    MUX21X1 U4392 (.IN1(next_mask_rr_arbiter31[j_rr_arbiter31[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter31), .Q(next_mask_rr_arbiter31[j_rr_arbiter31[0]]));
    MUX21X1 U4393 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U4394 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b1), .S(secondif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));
    NAND2X1 U4395 ( .IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(_sv2v_jump_rr_rr_arbiter31[1]), .QN(fourthif_rr_arbiter31) );
    MUX21X1 U4396 (.IN1(_sv2v_jump_rr_rr_arbiter31[0]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[0]));
    MUX21X1 U4397 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(fourthif_rr_arbiter31), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    MUX21X1 U4398 (.IN1(_sv2v_jump_rr_rr_arbiter31[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter31[1]));

    DFFX2 U4399 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter31) );
    DFFX2 U4400 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter31) );
    MUX21X1 U4401 (.IN1(mask_ff_rr_arbiter31[0]), .IN2(next_mask_rr_arbiter31[0]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[0]));
    MUX21X1 U4402 (.IN1(mask_ff_rr_arbiter31[1]), .IN2(next_mask_rr_arbiter31[1]), .S(tail_flit_im_output_module3[1]), .Q(temp_mask_ff_rr_arbiter3311[1]));
    MUX21X1 U4403 (.IN1(temp_mask_ff_rr_arbiter3311), .IN2(1'sb1), .S(arst_value_rr_arbiter31), .Q(mask_ff_rr_arbiter31[0]));





    BUFX1 U4404 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[0]) );
    BUFX1 U4405 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter132[1]) );
    BUFX1 U4406 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4407 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4408 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    XNOR2X1 U4409 ( .IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter132) );
    MUX21X1 U4410 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U4411 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    INVX1 U4412 ( .A(i_high_prior_arbiter132[0]), .Y(i_0_not_high_prior_arbiter132) );
    MUX21X1 U4413 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter132), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[0]);
    MUX21X1 U4414 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter132[0]), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(raw_grant[1]);
    MUX21X1 U4415 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U4416 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b1), .S(valid_from_im_output_module3[11:8][i_high_prior_arbiter132[0]]), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    NAND2X1 U4417 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(_sv2v_jump_high_prior_arbiter132[1]), .QN(nandres_high_prior_arbiter132) );
    MUX21X1 U4418 (.IN1(_sv2v_jump_high_prior_arbiter132[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[0]));
    MUX21X1 U4419 (.IN1(_sv2v_jump_high_prior_arbiter132[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter132), .Q(_sv2v_jump_high_prior_arbiter132[1]));
    HADDX1 U4420 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U4421 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );
    HADDX1 U4422 ( .A0(i_high_prior_arbiter132[0]), .B0(1'b1), .C1(i_high_prior_arbiter132[1]), .SO(i_high_prior_arbiter132[0]) );



    BUFX1 U4423 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[0]) );
    BUFX1 U4424 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter232[1]) );
    BUFX1 U4425 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4426 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4427 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    XNOR2X1 U4428 ( .IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter232) );
    MUX21X1 U4429 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U4430 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    INVX1 U4431 ( .A(i_high_prior_arbiter232[0]), .Y(i_0_not_high_prior_arbiter232) );
    MUX21X1 U4432 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter232), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[0]);
    MUX21X1 U4433 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter232[0]), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(masked_grant[1]);
    MUX21X1 U4434 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U4435 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter232[0]]), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    NAND2X1 U4436 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(_sv2v_jump_high_prior_arbiter232[1]), .QN(nandres_high_prior_arbiter232) );
    MUX21X1 U4437 (.IN1(_sv2v_jump_high_prior_arbiter232[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[0]));
    MUX21X1 U4438 (.IN1(_sv2v_jump_high_prior_arbiter232[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter232), .Q(_sv2v_jump_high_prior_arbiter232[1]));
    HADDX1 U4439 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U4440 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    HADDX1 U4441 ( .A0(i_high_prior_arbiter232[0]), .B0(1'b1), .C1(i_high_prior_arbiter232[1]), .SO(i_high_prior_arbiter232[0]) );
    

    BUFX1 U4442 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[0]) );
    BUFX1 U4443 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter32[1]) );
    AND2X1 U4444 ( .A(mask_ff_rr_arbiter32[0]), .B(valid_from_im_output_module3[11:8][0]), .Y(mask_req_rr_arbiter32[0]) );
    AND2X1 U4445 ( .A(mask_ff_rr_arbiter32[1]), .B(valid_from_im_output_module3[11:8][1]), .Y(mask_req_rr_arbiter32[1]) );
    BUFX1 U4446 ( .A(mask_ff_rr_arbiter32[0]), .Y(next_mask_rr_arbiter32[0]) );
    BUFX1 U4447 ( .A(mask_ff_rr_arbiter32[1]), .Y(next_mask_rr_arbiter32[1]) );
    XNOR2X1 U4448 ( .IN1(mask_req_rr_arbiter32[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter32) );
    XNOR2X1 U4449 ( .IN1(mask_req_rr_arbiter32[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter32) );
    MUX21X1 U4450 (.IN1(masked_grant_rr_arbiter32[0]), .IN2(raw_grant_rr_arbiter32[0]), .S(xnor0res_rr_arbiter32), .Q(grant_im_output_module3[11:8][0]));
    MUX21X1 U4451 (.IN1(masked_grant_rr_arbiter32[1]), .IN2(raw_grant_rr_arbiter32[1]), .S(xnor1res_rr_arbiter32), .Q(grant_im_output_module3[11:8][1]));

    BUFX1 U4452 ( .A(1'b0), .Y(i_rr_arbiter32[1]) );
    MUX21X1 U4453 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter32[0]));

    AND2X1 U4454 ( .A(_sv2v_jump_rr_rr_arbiter32[1]), .B(1'b0), .Y(firstif_rr_arbiter32) );
    MUX21X1 U4455 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U4456 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(firstif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    AND2X1 U4457 ( .A(firstif_rr_arbiter32), .B(grant_im_output_module3[11:8][i_rr_arbiter32[0]]), .Y(secondif_rr_arbiter32) );
    MUX21X1 U4458 (.IN1(next_mask_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[0]));
    MUX21X1 U4459 (.IN1(next_mask_rr_arbiter32[1]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(next_mask_rr_arbiter32[1]));
    MUX21X1 U4460 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter32[0]), .Q(j_rr_arbiter32[0]));
    AND2X1 U4461 ( .A(secondif_rr_arbiter32), .B(j_rr_arbiter32[0]), .Y(thirdif_rr_arbiter32) );
    MUX21X1 U4462 (.IN1(next_mask_rr_arbiter32[j_rr_arbiter32[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter32), .Q(next_mask_rr_arbiter32[j_rr_arbiter32[0]]));
    MUX21X1 U4463 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U4464 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b1), .S(secondif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));
    NAND2X1 U4465 ( .IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(_sv2v_jump_rr_rr_arbiter32[1]), .QN(fourthif_rr_arbiter32) );
    MUX21X1 U4466 (.IN1(_sv2v_jump_rr_rr_arbiter32[0]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[0]));
    MUX21X1 U4467 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(fourthif_rr_arbiter32), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    MUX21X1 U4468 (.IN1(_sv2v_jump_rr_rr_arbiter32[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter32[1]));

    DFFX2 U4469 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter32) );
    DFFX2 U4470 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter32) );
    MUX21X1 U4471 (.IN1(mask_ff_rr_arbiter32[0]), .IN2(next_mask_rr_arbiter32[0]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[0]));
    MUX21X1 U4472 (.IN1(mask_ff_rr_arbiter32[1]), .IN2(next_mask_rr_arbiter32[1]), .S(tail_flit_im_output_module3[2]), .Q(temp_mask_ff_rr_arbiter3322[1]));
    MUX21X1 U4473 (.IN1(temp_mask_ff_rr_arbiter3322), .IN2(1'sb1), .S(arst_value_rr_arbiter32), .Q(mask_ff_rr_arbiter32[0]));


    XNOR2X1 U4474 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37]), .IN2(vc_channel_output_module3[1]), .QN(xnor1resu1_output_module3) );
    XNOR2X1 U4475 ( .IN1(int_map_req_v[480:444][in_mod_output_module3[1:0]*37-1]), .IN2(vc_channel_output_module3[0]), .QN(xnor2resu1_output_module3) );
    AND2X1 U4476 ( .IN1(xnor1resu1_output_module3), .IN2(xnor2resu1_output_module3), .Q(and1resu1_output_module3) );
    MUX21X1 U4477 (.IN1(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]), .IN2(1'b1), .S(and1resu1_output_module3), .Q(valid_from_im_output_module3[(vc_channel_output_module3[1:0]*4) + in_mod_output_module3[1:0]]);
    HADDX1 U4478 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4479 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4480 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4481 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4482 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4483 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4484 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4485 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4486 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4487 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );  
    HADDX1 U4488 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4489 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4490 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4491 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) ); 
    XOR2X1 U4492 ( .IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .Q(xor1resu1_output_module3) );
    MUX21X1 U4493 (.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[0]));
    MUX21X1 U4494 (.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3[1]));
    MUX21X1 U4495 (.IN1(_sv2v_jump_output_module3_1[0]), .IN2(_sv2v_jump_output_module3[0]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[0]));
    MUX21X1 U4496 (.IN1(_sv2v_jump_output_module3_1[1]), .IN2(_sv2v_jump_output_module3[1]), .S(xor1resu1_output_module3), .Q(_sv2v_jump_output_module3_1[1]));
    AND2X1 U4497 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[vc_channel_output_module3[1:0]*4+in_mod_output_module3[1:0]]), .Q(and2resu1_output_module3) );

    MUX21X1 U4498(.IN1(head_flit_output_module3[3]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+3]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[3]));
    MUX21X1 U4499(.IN1(head_flit_output_module3[4]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+4]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[4]));
    MUX21X1 U4500(.IN1(head_flit_output_module3[5]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+5]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[5]));
    MUX21X1 U4501(.IN1(head_flit_output_module3[6]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+6]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[6]));
    MUX21X1 U4502(.IN1(head_flit_output_module3[7]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+7]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[7]));
    MUX21X1 U4503(.IN1(head_flit_output_module3[8]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+8]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[8]));
    MUX21X1 U4504(.IN1(head_flit_output_module3[9]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+9]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[9]));
    MUX21X1 U4505(.IN1(head_flit_output_module3[10]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+10]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[10]));
    MUX21X1 U4506(.IN1(head_flit_output_module3[11]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+11]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[11]));
    MUX21X1 U4507(.IN1(head_flit_output_module3[12]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+12]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[12]));
    MUX21X1 U4508(.IN1(head_flit_output_module3[13]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+13]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[13]));
    MUX21X1 U4509(.IN1(head_flit_output_module3[14]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+14]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[14]));
    MUX21X1 U4510(.IN1(head_flit_output_module3[15]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+15]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[15]));
    MUX21X1 U4511(.IN1(head_flit_output_module3[16]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+16]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[16]));
    MUX21X1 U4512(.IN1(head_flit_output_module3[17]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+17]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[17]));
    MUX21X1 U4513(.IN1(head_flit_output_module3[18]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+18]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[18]));
    MUX21X1 U4514(.IN1(head_flit_output_module3[19]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+19]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[19]));
    MUX21X1 U4515(.IN1(head_flit_output_module3[20]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+20]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[20]));
    MUX21X1 U4516(.IN1(head_flit_output_module3[21]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+21]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[21]));
    MUX21X1 U4517(.IN1(head_flit_output_module3[22]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+22]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[22]));
    MUX21X1 U4518(.IN1(head_flit_output_module3[23]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+23]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[23]));
    MUX21X1 U4519(.IN1(head_flit_output_module3[24]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+24]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[24]));
    MUX21X1 U4520(.IN1(head_flit_output_module3[25]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+25]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[25]));
    MUX21X1 U4521(.IN1(head_flit_output_module3[26]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+26]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[26]));
    MUX21X1 U4522(.IN1(head_flit_output_module3[27]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+27]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[27]));
    MUX21X1 U4523(.IN1(head_flit_output_module3[28]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+28]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[28]));
    MUX21X1 U4524(.IN1(head_flit_output_module3[29]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+29]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[29]));
    MUX21X1 U4525(.IN1(head_flit_output_module3[30]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+30]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[30]));
    MUX21X1 U4526(.IN1(head_flit_output_module3[31]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+31]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[31]));
    MUX21X1 U4527(.IN1(head_flit_output_module3[32]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+32]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[32]));
    MUX21X1 U4528(.IN1(head_flit_output_module3[33]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+33]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[33]));
    MUX21X1 U4529(.IN1(head_flit_output_module3[34]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+34]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[34]));
    MUX21X1 U4530(.IN1(head_flit_output_module3[35]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+35]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[35]));
    MUX21X1 U4531(.IN1(head_flit_output_module3[36]), .IN2(int_map_req_v[480:444][in_mod_output_module3[1:0]*37+36]), .S(and2resu1_output_module3) ,.Q(head_flit_output_module3[36]));

    INVX1 U4532 ( .A(head_flit_output_module3[32]), .Y(head_flit_output_module3_32_not_output_module3) );
    AND2X1 U4533 ( .IN1(head_flit_output_module3_32_not_output_module3), .IN2(head_flit_output_module3[33]), .Q(and3resu1_output_module3) );
    NOR4X1 U4534 (.IN1(head_flit_output_module3[29]), .IN2(head_flit_output_module3[28]), .IN3(head_flit_output_module3[27]), .IN4(head_flit_output_module3[26]), .Q(nor23resu1_output_module3) );
    NOR4X1 U4535 (.IN1(head_flit_output_module3[25]), .IN2(head_flit_output_module3[24]), .IN3(head_flit_output_module3[23]), .IN4(head_flit_output_module3[22]), .Q(nor23resu2_output_module3) );
    AND2X1 U4536 ( .IN1(nor23resu1_output_module3), .IN2(nor23resu2_output_module3), .Q(and4resu1_output_module3) );
    NOR2X1 U4537 (.IN1(head_flit_output_module3[33]), .IN2(head_flit_output_module3[32]), .Q(nor23resu3_output_module3) );
    AND2X1 U4538 ( .IN1(nor23resu3_output_module3), .IN2(and4resu1_output_module3), .Q(and5resu1_output_module3) );    
    OR2X1 U4539 (.IN1(and3resu1_output_module3), .IN2(nor23resu3_output_module3), .Q(or12resu12_output_module3) );
    AND2X1 U4540 ( .IN1(ext_resp_v_i[4:3][0]), .IN2(or12resu12_output_module3), .Q(and6resu1_output_module3) );    
    MUX21X1 U4541(.IN1(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]), .IN2(and6resu1_output_module3), .S(and2resu1_output_module3) ,.Q(tail_flit_im_output_module3[vc_channel_output_module3[1:0]]);
    MUX21X1 U4542(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4543(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and2resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    NAND2X1 U4544(.A(_sv2v_jump_output_module3[0]),.B(_sv2v_jump_output_module3[1]),.Y(nand1resu_output_module3));

    AND2X1 U4545 ( .IN1(xor1resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and7resu1) );    
    MUX21X1 U4546(.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4547(.IN1(_sv2v_jump_output_module3[1]), .IN2(_sv2v_jump_output_module3_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    MUX21X1 U4548(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4549(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module3[1]);

    HADDX1 U4550 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4551 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4552 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4553 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4554 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4555 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4556 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4557 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4558 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4559 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4560 ( .A0(vc_channel_output_module3[0]), .B0(1'b1), .C1(vc_channel_output_module3[1]), .SO(vc_channel_output_module3[0]) );
    HADDX1 U4561 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4562 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4563 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );
    HADDX1 U4564 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(in_mod_output_module3[1]), .SO(in_mod_output_module3[0]) );



    BUFX1 U4565(.A(1'b0), .Y(_sv2v_jump_output_module3[0]));
    BUFX1 U4566(.A(1'b0), .Y(_sv2v_jump_output_module3[1]));
    AND2X1 U4567 ( .IN1(xor1resu1_output_module3), .IN2(grant_im_output_module3[i_output_module3[1:0] * 4+:4]), .Q(and8resu1_output_module3) );    
    MUX21X1 U4568(.IN1(vc_ch_act_out_output_module3[0]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[0]);
    MUX21X1 U4569(.IN1(vc_ch_act_out_output_module3[1]), .IN2(i_output_module3[1:0]), .S(and8resu1_output_module3) ,.Q(vc_ch_act_out_output_module3[1]);
    MUX21X1 U4570(.IN1(req_out_output_module3), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(req_out_output_module3);
    MUX21X1 U4571(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4572(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and8resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);
    HADDX1 U4573 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U4574 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    HADDX1 U4575 ( .A0(in_mod_output_module3[0]), .B0(1'b1), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );

    NOR2X1 U4576 (.IN1(_sv2v_jump_output_module3[0]), .IN2(_sv2v_jump_output_module3[1]), .Q(norfinresu1_output_module3) );
    AND2X1 U4577 ( .IN1(norfinresu1_output_module3), .IN2(req_out_output_module3), .Q(and9resu1_output_module3) );    
    HADDX1 U4578 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module3[1]), .SO(i_output_module3[0]) );
    AND2X1 U4579 ( .IN1(and9resu1_output_module3), .IN2(grant_im_output_module3[(vc_ch_act_out_output_module3 * 4) + i_output_module3[1:0]]), .Q(and10resu1_output_module3) );    

    MUX21X1 U4580(.IN1(ext_req_v_o[147:111][3]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+3]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][3]));
    MUX21X1 U4581(.IN1(ext_req_v_o[147:111][4]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+4]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][4]));
    MUX21X1 U4582(.IN1(ext_req_v_o[147:111][5]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+5]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][5]));
    MUX21X1 U4583(.IN1(ext_req_v_o[147:111][6]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+6]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][6]));
    MUX21X1 U4584(.IN1(ext_req_v_o[147:111][7]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+7]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][7]));
    MUX21X1 U4585(.IN1(ext_req_v_o[147:111][8]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+8]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][8]));
    MUX21X1 U4586(.IN1(ext_req_v_o[147:111][9]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+9]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][9]));
    MUX21X1 U4587(.IN1(ext_req_v_o[147:111][10]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+10]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][10]));
    MUX21X1 U4588(.IN1(ext_req_v_o[147:111][11]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+11]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][11]));
    MUX21X1 U4589(.IN1(ext_req_v_o[147:111][12]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+12]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][12]));
    MUX21X1 U4590(.IN1(ext_req_v_o[147:111][13]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+13]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][13]));
    MUX21X1 U4591(.IN1(ext_req_v_o[147:111][14]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+14]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][14]));
    MUX21X1 U4592(.IN1(ext_req_v_o[147:111][15]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+15]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][15]));
    MUX21X1 U4593(.IN1(ext_req_v_o[147:111][16]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+16]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][16]));
    MUX21X1 U4594(.IN1(ext_req_v_o[147:111][17]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+17]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][17]));
    MUX21X1 U4595(.IN1(ext_req_v_o[147:111][18]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+18]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][18]));
    MUX21X1 U4596(.IN1(ext_req_v_o[147:111][19]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+19]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][19]));
    MUX21X1 U4597(.IN1(ext_req_v_o[147:111][20]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+20]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][20]));
    MUX21X1 U4598(.IN1(ext_req_v_o[147:111][21]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+21]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][21]));
    MUX21X1 U4599(.IN1(ext_req_v_o[147:111][22]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+22]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][22]));
    MUX21X1 U4600(.IN1(ext_req_v_o[147:111][23]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+23]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][23]));
    MUX21X1 U4601(.IN1(ext_req_v_o[147:111][24]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+24]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][24]));
    MUX21X1 U4602(.IN1(ext_req_v_o[147:111][25]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+25]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][25]));
    MUX21X1 U4603(.IN1(ext_req_v_o[147:111][26]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+26]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][26]));
    MUX21X1 U4604(.IN1(ext_req_v_o[147:111][27]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+27]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][27]));
    MUX21X1 U4605(.IN1(ext_req_v_o[147:111][28]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+28]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][28]));
    MUX21X1 U4606(.IN1(ext_req_v_o[147:111][29]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+29]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][29]));
    MUX21X1 U4607(.IN1(ext_req_v_o[147:111][30]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+30]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][30]));
    MUX21X1 U4608(.IN1(ext_req_v_o[147:111][31]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+31]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][31]));
    MUX21X1 U4609(.IN1(ext_req_v_o[147:111][32]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+32]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][32]));
    MUX21X1 U4610(.IN1(ext_req_v_o[147:111][33]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+33]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][33]));
    MUX21X1 U4611(.IN1(ext_req_v_o[147:111][34]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+34]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][34]));
    MUX21X1 U4612(.IN1(ext_req_v_o[147:111][35]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+35]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][35]));
    MUX21X1 U4613(.IN1(ext_req_v_o[147:111][36]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37+36]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][36]));

    MUX21X1 U4614(.IN1(ext_req_v_o[147:111][0]), .IN2(int_map_req_v[480:444][i_output_module3[1:0]*37]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][0]);
    MUX21X1 U4615(.IN1(ext_req_v_o[147:111][1]), .IN2(vc_ch_act_out_output_module3[0]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][1]);
    MUX21X1 U4616(.IN1(ext_req_v_o[147:111][2]), .IN2(vc_ch_act_out_output_module3[1]), .S(and10resu1_output_module3) ,.Q(ext_req_v_o[147:111][2]);    
    MUX21X1 U4617(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4618(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b1), .S(and10resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    

    AND2X1 U4619 ( .IN1(and9resu1_output_module3), .IN2(nand1resu_output_module3), .Q(and11resu1_output_module3) );    
    MUX21X1 U4620(.IN1(_sv2v_jump_output_module3[0]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[0]);
    MUX21X1 U4621(.IN1(_sv2v_jump_output_module3[1]), .IN2(1'b0), .S(and11resu1_output_module3) ,.Q(_sv2v_jump_output_module3[1]);    







    BUFX1 U4622 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[0]) );
    BUFX1 U4623 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter14[1]) );
    BUFX1 U4624 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4625 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4626 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    XNOR2X1 U4627 ( .IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter14) );
    MUX21X1 U4628 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U4629 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    INVX1 U4630 ( .A(i_high_prior_arbiter14[0]), .Y(i_0_not_high_prior_arbiter14) );
    MUX21X1 U4631 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter14), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[0]);
    MUX21X1 U4632 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter14[0]), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(raw_grant[1]);
    MUX21X1 U4633 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U4634 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b1), .S(valid_from_im_output_module4[3:0][i_high_prior_arbiter14[0]]), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    NAND2X1 U4635 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(_sv2v_jump_high_prior_arbiter14[1]), .QN(nandres_high_prior_arbiter14) );
    MUX21X1 U4636 (.IN1(_sv2v_jump_high_prior_arbiter14[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[0]));
    MUX21X1 U4637 (.IN1(_sv2v_jump_high_prior_arbiter14[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter14), .Q(_sv2v_jump_high_prior_arbiter14[1]));
    HADDX1 U4638 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U4639 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );
    HADDX1 U4640 ( .A0(i_high_prior_arbiter14[0]), .B0(1'b1), .C1(i_high_prior_arbiter14[1]), .SO(i_high_prior_arbiter14[0]) );



    BUFX1 U4641 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[0]) );
    BUFX1 U4642 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter24[1]) );
    BUFX1 U4643 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4644 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4645 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    XNOR2X1 U4646 ( .IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter24) );
    MUX21X1 U4647 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U4648 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    INVX1 U4649 ( .A(i_high_prior_arbiter24[0]), .Y(i_0_not_high_prior_arbiter24) );
    MUX21X1 U4650 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter24), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[0]);
    MUX21X1 U4651 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter24[0]), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(masked_grant[1]);
    MUX21X1 U4652 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U4653 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter24[0]]), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    NAND2X1 U4654 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(_sv2v_jump_high_prior_arbiter24[1]), .QN(nandres_high_prior_arbiter24) );
    MUX21X1 U4655 (.IN1(_sv2v_jump_high_prior_arbiter24[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[0]));
    MUX21X1 U4656 (.IN1(_sv2v_jump_high_prior_arbiter24[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter24), .Q(_sv2v_jump_high_prior_arbiter24[1]));
    HADDX1 U4657 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U4658 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    HADDX1 U4659 ( .A0(i_high_prior_arbiter24[0]), .B0(1'b1), .C1(i_high_prior_arbiter24[1]), .SO(i_high_prior_arbiter24[0]) );
    

    BUFX1 U4660 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[0]) );
    BUFX1 U4661 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter4[1]) );
    AND2X1 U4662 ( .A(mask_ff_rr_arbiter4[0]), .B(valid_from_im_output_module4[3:0][0]), .Y(mask_req_rr_arbiter4[0]) );
    AND2X1 U4663 ( .A(mask_ff_rr_arbiter4[1]), .B(valid_from_im_output_module4[3:0][1]), .Y(mask_req_rr_arbiter4[1]) );
    BUFX1 U4664 ( .A(mask_ff_rr_arbiter4[0]), .Y(next_mask_rr_arbiter4[0]) );
    BUFX1 U4665 ( .A(mask_ff_rr_arbiter4[1]), .Y(next_mask_rr_arbiter4[1]) );
    XNOR2X1 U4666 ( .IN1(mask_req_rr_arbiter4[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter4) );
    XNOR2X1 U4667 ( .IN1(mask_req_rr_arbiter4[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter4) );
    MUX21X1 U4668 (.IN1(masked_grant_rr_arbiter4[0]), .IN2(raw_grant_rr_arbiter4[0]), .S(xnor0res_rr_arbiter4), .Q(grant_im_output_module4[3:0][0]));
    MUX21X1 U4669 (.IN1(masked_grant_rr_arbiter4[1]), .IN2(raw_grant_rr_arbiter4[1]), .S(xnor1res_rr_arbiter4), .Q(grant_im_output_module4[3:0][1]));

    BUFX1 U4670 ( .A(1'b0), .Y(i_rr_arbiter4[1]) );
    MUX21X1 U4671 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter4[0]));

    AND2X1 U4672 ( .A(_sv2v_jump_rr_rr_arbiter4[1]), .B(1'b0), .Y(firstif_rr_arbiter4) );
    MUX21X1 U4673 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U4674 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(firstif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    AND2X1 U4675 ( .A(firstif_rr_arbiter4), .B(grant_im_output_module4[3:0][i_rr_arbiter4[0]]), .Y(secondif_rr_arbiter4) );
    MUX21X1 U4676 (.IN1(next_mask_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[0]));
    MUX21X1 U4677 (.IN1(next_mask_rr_arbiter4[1]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(next_mask_rr_arbiter4[1]));
    MUX21X1 U4678 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter4[0]), .Q(j_rr_arbiter4[0]));
    AND2X1 U4679 ( .A(secondif_rr_arbiter4), .B(j_rr_arbiter4[0]), .Y(thirdif_rr_arbiter4) );
    MUX21X1 U4680 (.IN1(next_mask_rr_arbiter4[j_rr_arbiter4[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter4), .Q(next_mask_rr_arbiter4[j_rr_arbiter4[0]]));
    MUX21X1 U4681 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U4682 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b1), .S(secondif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));
    NAND2X1 U4683 ( .IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(_sv2v_jump_rr_rr_arbiter4[1]), .QN(fourthif_rr_arbiter4) );
    MUX21X1 U4684 (.IN1(_sv2v_jump_rr_rr_arbiter4[0]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[0]));
    MUX21X1 U4685 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(fourthif_rr_arbiter4), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    MUX21X1 U4686 (.IN1(_sv2v_jump_rr_rr_arbiter4[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter4[1]));

    DFFX2 U4687 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter4) );
    DFFX2 U4688 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter4) );
    MUX21X1 U4689 (.IN1(mask_ff_rr_arbiter4[0]), .IN2(next_mask_rr_arbiter4[0]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[0]));
    MUX21X1 U4690 (.IN1(mask_ff_rr_arbiter4[1]), .IN2(next_mask_rr_arbiter4[1]), .S(tail_flit_im_output_module4[0]), .Q(temp_mask_ff_rr_arbiter44[1]));
    MUX21X1 U4691 (.IN1(temp_mask_ff_rr_arbiter44), .IN2(1'sb1), .S(arst_value_rr_arbiter4), .Q(mask_ff_rr_arbiter4[0]));



    BUFX1 U4692 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[0]) );
    BUFX1 U4693 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter141[1]) );
    BUFX1 U4694 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4695 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4696 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    XNOR2X1 U4697 ( .IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter141) );
    MUX21X1 U4698 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U4699 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    INVX1 U4700 ( .A(i_high_prior_arbiter141[0]), .Y(i_0_not_high_prior_arbiter141) );
    MUX21X1 U4701 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter141), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[0]);
    MUX21X1 U4702 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter141[0]), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(raw_grant[1]);
    MUX21X1 U4703 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U4704 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b1), .S(valid_from_im_output_module4[7:4][i_high_prior_arbiter141[0]]), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    NAND2X1 U4705 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(_sv2v_jump_high_prior_arbiter141[1]), .QN(nandres_high_prior_arbiter141) );
    MUX21X1 U4706 (.IN1(_sv2v_jump_high_prior_arbiter141[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[0]));
    MUX21X1 U4707 (.IN1(_sv2v_jump_high_prior_arbiter141[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter141), .Q(_sv2v_jump_high_prior_arbiter141[1]));
    HADDX1 U4708 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U4709 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );
    HADDX1 U4710 ( .A0(i_high_prior_arbiter141[0]), .B0(1'b1), .C1(i_high_prior_arbiter141[1]), .SO(i_high_prior_arbiter141[0]) );



    BUFX1 U4711 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[0]) );
    BUFX1 U4712 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter241[1]) );
    BUFX1 U4713 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4714 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4715 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    XNOR2X1 U4716 ( .IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter2414) );
    MUX21X1 U4717 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U4718 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    INVX1 U4719 ( .A(i_high_prior_arbiter241[0]), .Y(i_0_not_high_prior_arbiter2414) );
    MUX21X1 U4720 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter2414), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[0]);
    MUX21X1 U4721 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter241[0]), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(masked_grant[1]);
    MUX21X1 U4722 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U4723 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter241[0]]), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    NAND2X1 U4724 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(_sv2v_jump_high_prior_arbiter241[1]), .QN(nandres_high_prior_arbiter2414) );
    MUX21X1 U4725 (.IN1(_sv2v_jump_high_prior_arbiter241[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[0]));
    MUX21X1 U4726 (.IN1(_sv2v_jump_high_prior_arbiter241[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter2414), .Q(_sv2v_jump_high_prior_arbiter241[1]));
    HADDX1 U4727 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U4728 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    HADDX1 U4729 ( .A0(i_high_prior_arbiter241[0]), .B0(1'b1), .C1(i_high_prior_arbiter241[1]), .SO(i_high_prior_arbiter241[0]) );
    

    BUFX1 U4730 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[0]) );
    BUFX1 U4731 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter41[1]) );
    AND2X1 U4732 ( .A(mask_ff_rr_arbiter41[0]), .B(valid_from_im_output_module4[7:4][0]), .Y(mask_req_rr_arbiter41[0]) );
    AND2X1 U4733 ( .A(mask_ff_rr_arbiter41[1]), .B(valid_from_im_output_module4[7:4][1]), .Y(mask_req_rr_arbiter41[1]) );
    BUFX1 U4734 ( .A(mask_ff_rr_arbiter41[0]), .Y(next_mask_rr_arbiter41[0]) );
    BUFX1 U4735 ( .A(mask_ff_rr_arbiter41[1]), .Y(next_mask_rr_arbiter41[1]) );
    XNOR2X1 U4736 ( .IN1(mask_req_rr_arbiter41[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter41) );
    XNOR2X1 U4737 ( .IN1(mask_req_rr_arbiter41[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter41) );
    MUX21X1 U4738 (.IN1(masked_grant_rr_arbiter41[0]), .IN2(raw_grant_rr_arbiter41[0]), .S(xnor0res_rr_arbiter41), .Q(grant_im_output_module4[7:4][0]));
    MUX21X1 U4739 (.IN1(masked_grant_rr_arbiter41[1]), .IN2(raw_grant_rr_arbiter41[1]), .S(xnor1res_rr_arbiter41), .Q(grant_im_output_module4[7:4][1]));

    BUFX1 U4740 ( .A(1'b0), .Y(i_rr_arbiter41[1]) );
    MUX21X1 U4741 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter41[0]));

    AND2X1 U4742 ( .A(_sv2v_jump_rr_rr_arbiter41[1]), .B(1'b0), .Y(firstif_rr_arbiter41) );
    MUX21X1 U4743 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U4744 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(firstif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    AND2X1 U4745 ( .A(firstif_rr_arbiter41), .B(grant_im_output_module4[7:4][i_rr_arbiter41[0]]), .Y(secondif_rr_arbiter41) );
    MUX21X1 U4746 (.IN1(next_mask_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[0]));
    MUX21X1 U4747 (.IN1(next_mask_rr_arbiter41[1]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(next_mask_rr_arbiter41[1]));
    MUX21X1 U4748 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter41[0]), .Q(j_rr_arbiter41[0]));
    AND2X1 U4749 ( .A(secondif_rr_arbiter41), .B(j_rr_arbiter41[0]), .Y(thirdif_rr_arbiter41) );
    MUX21X1 U4750 (.IN1(next_mask_rr_arbiter41[j_rr_arbiter41[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter41), .Q(next_mask_rr_arbiter41[j_rr_arbiter41[0]]));
    MUX21X1 U4751 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U4752 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b1), .S(secondif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));
    NAND2X1 U4753 ( .IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(_sv2v_jump_rr_rr_arbiter41[1]), .QN(fourthif_rr_arbiter41) );
    MUX21X1 U4754 (.IN1(_sv2v_jump_rr_rr_arbiter41[0]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[0]));
    MUX21X1 U4755 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(fourthif_rr_arbiter41), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    MUX21X1 U4756 (.IN1(_sv2v_jump_rr_rr_arbiter41[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter41[1]));

    DFFX2 U4757 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter41) );
    DFFX2 U4758 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter41) );
    MUX21X1 U4759 (.IN1(mask_ff_rr_arbiter41[0]), .IN2(next_mask_rr_arbiter41[0]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[0]));
    MUX21X1 U4760 (.IN1(mask_ff_rr_arbiter41[1]), .IN2(next_mask_rr_arbiter41[1]), .S(tail_flit_im_output_module4[1]), .Q(temp_mask_ff_rr_arbiter4411[1]));
    MUX21X1 U4761 (.IN1(temp_mask_ff_rr_arbiter4411), .IN2(1'sb1), .S(arst_value_rr_arbiter41), .Q(mask_ff_rr_arbiter41[0]));





    BUFX1 U4762 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[0]) );
    BUFX1 U4763 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter142[1]) );
    BUFX1 U4764 ( .A(1'b0), .Y(raw_grant[0]) );
    BUFX1 U4765 ( .A(1'b0), .Y(raw_grant[1]) );
    HADDX1 U4766 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    XNOR2X1 U4767 ( .IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter142) );
    MUX21X1 U4768 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U4769 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    INVX1 U4770 ( .A(i_high_prior_arbiter142[0]), .Y(i_0_not_high_prior_arbiter142) );
    MUX21X1 U4771 (.IN1(raw_grant[0]), .IN2(i_0_not_high_prior_arbiter142), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[0]);
    MUX21X1 U4772 (.IN1(raw_grant[1]), .IN2(i_high_prior_arbiter142[0]), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(raw_grant[1]);
    MUX21X1 U4773 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U4774 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b1), .S(valid_from_im_output_module4[11:8][i_high_prior_arbiter142[0]]), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    NAND2X1 U4775 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(_sv2v_jump_high_prior_arbiter142[1]), .QN(nandres_high_prior_arbiter142) );
    MUX21X1 U4776 (.IN1(_sv2v_jump_high_prior_arbiter142[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[0]));
    MUX21X1 U4777 (.IN1(_sv2v_jump_high_prior_arbiter142[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter142), .Q(_sv2v_jump_high_prior_arbiter142[1]));
    HADDX1 U4778 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U4779 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );
    HADDX1 U4780 ( .A0(i_high_prior_arbiter142[0]), .B0(1'b1), .C1(i_high_prior_arbiter142[1]), .SO(i_high_prior_arbiter142[0]) );



    BUFX1 U4781 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[0]) );
    BUFX1 U4782 ( .A(1'b0), .Y(_sv2v_jump_high_prior_arbiter242[1]) );
    BUFX1 U4783 ( .A(1'b0), .Y(masked_grant[0]) );
    BUFX1 U4784 ( .A(1'b0), .Y(masked_grant[1]) );
    HADDX1 U4785 ( .A0(1'b0), .B0(1'b0), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    XNOR2X1 U4786 ( .IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .Q(xnores_high_prior_arbiter242) );
    MUX21X1 U4787 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U4788 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(xnores_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    INVX1 U4789 ( .A(i_high_prior_arbiter242[0]), .Y(i_0_not_high_prior_arbiter242) );
    MUX21X1 U4790 (.IN1(masked_grant[0]), .IN2(i_0_not_high_prior_arbiter242), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[0]);
    MUX21X1 U4791 (.IN1(masked_grant[1]), .IN2(i_high_prior_arbiter242[0]), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(masked_grant[1]);
    MUX21X1 U4792 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U4793 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b1), .S(mask_req[i_high_prior_arbiter242[0]]), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    NAND2X1 U4794 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(_sv2v_jump_high_prior_arbiter242[1]), .QN(nandres_high_prior_arbiter242) );
    MUX21X1 U4795 (.IN1(_sv2v_jump_high_prior_arbiter242[0]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[0]));
    MUX21X1 U4796 (.IN1(_sv2v_jump_high_prior_arbiter242[1]), .IN2(1'b0), .S(nandres_high_prior_arbiter242), .Q(_sv2v_jump_high_prior_arbiter242[1]));
    HADDX1 U4797 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U4798 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    HADDX1 U4799 ( .A0(i_high_prior_arbiter242[0]), .B0(1'b1), .C1(i_high_prior_arbiter242[1]), .SO(i_high_prior_arbiter242[0]) );
    

    BUFX1 U4800 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[0]) );
    BUFX1 U4801 ( .A(1'b0), .Y(_sv2v_jump_rr_rr_arbiter42[1]) );
    AND2X1 U4802 ( .A(mask_ff_rr_arbiter42[0]), .B(valid_from_im_output_module4[11:8][0]), .Y(mask_req_rr_arbiter42[0]) );
    AND2X1 U4803 ( .A(mask_ff_rr_arbiter42[1]), .B(valid_from_im_output_module4[11:8][1]), .Y(mask_req_rr_arbiter42[1]) );
    BUFX1 U4804 ( .A(mask_ff_rr_arbiter42[0]), .Y(next_mask_rr_arbiter42[0]) );
    BUFX1 U4805 ( .A(mask_ff_rr_arbiter42[1]), .Y(next_mask_rr_arbiter42[1]) );
    XNOR2X1 U4806 ( .IN1(mask_req_rr_arbiter42[0]), .IN2(1'b0), .Q(xnor0res_rr_arbiter42) );
    XNOR2X1 U4807 ( .IN1(mask_req_rr_arbiter42[1]), .IN2(1'b0), .Q(xnor1res_rr_arbiter42) );
    MUX21X1 U4808 (.IN1(masked_grant_rr_arbiter42[0]), .IN2(raw_grant_rr_arbiter42[0]), .S(xnor0res_rr_arbiter42), .Q(grant_im_output_module4[11:8][0]));
    MUX21X1 U4809 (.IN1(masked_grant_rr_arbiter42[1]), .IN2(raw_grant_rr_arbiter42[1]), .S(xnor1res_rr_arbiter42), .Q(grant_im_output_module4[11:8][1]));

    BUFX1 U4810 ( .A(1'b0), .Y(i_rr_arbiter42[1]) );
    MUX21X1 U4811 (.IN1(1'b0), .IN2(1'b1), .S(clk), .Q(i_rr_arbiter42[0]));

    AND2X1 U4812 ( .A(_sv2v_jump_rr_rr_arbiter42[1]), .B(1'b0), .Y(firstif_rr_arbiter42) );
    MUX21X1 U4813 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U4814 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(firstif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    AND2X1 U4815 ( .A(firstif_rr_arbiter42), .B(grant_im_output_module4[11:8][i_rr_arbiter42[0]]), .Y(secondif_rr_arbiter42) );
    MUX21X1 U4816 (.IN1(next_mask_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[0]));
    MUX21X1 U4817 (.IN1(next_mask_rr_arbiter42[1]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(next_mask_rr_arbiter42[1]));
    MUX21X1 U4818 (.IN1(1'b1), .IN2(1'b0), .S(i_rr_arbiter42[0]), .Q(j_rr_arbiter42[0]));
    AND2X1 U4819 ( .A(secondif_rr_arbiter42), .B(j_rr_arbiter42[0]), .Y(thirdif_rr_arbiter42) );
    MUX21X1 U4820 (.IN1(next_mask_rr_arbiter42[j_rr_arbiter42[0]]), .IN2(1'b1), .S(thirdif_rr_arbiter42), .Q(next_mask_rr_arbiter42[j_rr_arbiter42[0]]));
    MUX21X1 U4821 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U4822 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b1), .S(secondif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));
    NAND2X1 U4823 ( .IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(_sv2v_jump_rr_rr_arbiter42[1]), .QN(fourthif_rr_arbiter42) );
    MUX21X1 U4824 (.IN1(_sv2v_jump_rr_rr_arbiter42[0]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[0]));
    MUX21X1 U4825 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(fourthif_rr_arbiter42), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    MUX21X1 U4826 (.IN1(_sv2v_jump_rr_rr_arbiter42[1]), .IN2(1'b0), .S(arst), .Q(_sv2v_jump_rr_rr_arbiter42[1]));

    DFFX2 U4827 ( .CLK(clk), .D(arst), .Q(arst_value_rr_arbiter42) );
    DFFX2 U4828 ( .CLK(arst), .D(arst), .Q(arst_value_rr_arbiter42) );
    MUX21X1 U4829 (.IN1(mask_ff_rr_arbiter42[0]), .IN2(next_mask_rr_arbiter42[0]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[0]));
    MUX21X1 U4830 (.IN1(mask_ff_rr_arbiter42[1]), .IN2(next_mask_rr_arbiter42[1]), .S(tail_flit_im_output_module4[2]), .Q(temp_mask_ff_rr_arbiter4422[1]));
    MUX21X1 U4831 (.IN1(temp_mask_ff_rr_arbiter4422), .IN2(1'sb1), .S(arst_value_rr_arbiter42), .Q(mask_ff_rr_arbiter42[0]));


    XNOR2X1 U4832 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37]), .IN2(vc_channel_output_module4[1]), .QN(xnor1resu1_output_module4) );
    XNOR2X1 U4833 ( .IN1(int_map_req_v[628:592][in_mod_output_module4[1:0]*37-1]), .IN2(vc_channel_output_module4[0]), .QN(xnor2resu1_output_module4) );
    AND2X1 U4834 ( .IN1(xnor1resu1_output_module4), .IN2(xnor2resu1_output_module4), .Q(and1resu1_output_module4) );
    MUX21X1 U4835 (.IN1(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]), .IN2(1'b1), .S(and1resu1_output_module4), .Q(valid_from_im_output_module4[(vc_channel_output_module4[1:0]*4) + in_mod_output_module4[1:0]]);
    HADDX1 U4836 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4837 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4838 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4839 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4840 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4841 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4842 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4843 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4844 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4845 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );  
    HADDX1 U4846 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4847 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4848 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4849 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) ); 
    XOR2X1 U4850 ( .IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .Q(xor1resu1_output_module4) );
    MUX21X1 U4851 (.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[0]));
    MUX21X1 U4852 (.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4[1]));
    MUX21X1 U4853 (.IN1(_sv2v_jump_output_module4_1[0]), .IN2(_sv2v_jump_output_module4[0]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[0]));
    MUX21X1 U4854 (.IN1(_sv2v_jump_output_module4_1[1]), .IN2(_sv2v_jump_output_module4[1]), .S(xor1resu1_output_module4), .Q(_sv2v_jump_output_module4_1[1]));
    AND2X1 U4855 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[vc_channel_output_module4[1:0]*4+in_mod_output_module4[1:0]]), .Q(and2resu1_output_module4) );

    MUX21X1 U4856(.IN1(head_flit_output_module4[3]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+3]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[3]));
    MUX21X1 U4857(.IN1(head_flit_output_module4[4]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+4]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[4]));
    MUX21X1 U4858(.IN1(head_flit_output_module4[5]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+5]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[5]));
    MUX21X1 U4859(.IN1(head_flit_output_module4[6]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+6]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[6]));
    MUX21X1 U4860(.IN1(head_flit_output_module4[7]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+7]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[7]));
    MUX21X1 U4861(.IN1(head_flit_output_module4[8]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+8]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[8]));
    MUX21X1 U4862(.IN1(head_flit_output_module4[9]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+9]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[9]));
    MUX21X1 U4863(.IN1(head_flit_output_module4[10]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+10]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[10]));
    MUX21X1 U4864(.IN1(head_flit_output_module4[11]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+11]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[11]));
    MUX21X1 U4865(.IN1(head_flit_output_module4[12]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+12]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[12]));
    MUX21X1 U4866(.IN1(head_flit_output_module4[13]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+13]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[13]));
    MUX21X1 U4867(.IN1(head_flit_output_module4[14]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+14]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[14]));
    MUX21X1 U4868(.IN1(head_flit_output_module4[15]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+15]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[15]));
    MUX21X1 U4869(.IN1(head_flit_output_module4[16]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+16]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[16]));
    MUX21X1 U4870(.IN1(head_flit_output_module4[17]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+17]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[17]));
    MUX21X1 U4871(.IN1(head_flit_output_module4[18]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+18]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[18]));
    MUX21X1 U4872(.IN1(head_flit_output_module4[19]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+19]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[19]));
    MUX21X1 U4873(.IN1(head_flit_output_module4[20]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+20]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[20]));
    MUX21X1 U4874(.IN1(head_flit_output_module4[21]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+21]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[21]));
    MUX21X1 U4875(.IN1(head_flit_output_module4[22]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+22]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[22]));
    MUX21X1 U4876(.IN1(head_flit_output_module4[23]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+23]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[23]));
    MUX21X1 U4877(.IN1(head_flit_output_module4[24]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+24]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[24]));
    MUX21X1 U4878(.IN1(head_flit_output_module4[25]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+25]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[25]));
    MUX21X1 U4879(.IN1(head_flit_output_module4[26]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+26]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[26]));
    MUX21X1 U4880(.IN1(head_flit_output_module4[27]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+27]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[27]));
    MUX21X1 U4881(.IN1(head_flit_output_module4[28]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+28]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[28]));
    MUX21X1 U4882(.IN1(head_flit_output_module4[29]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+29]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[29]));
    MUX21X1 U4883(.IN1(head_flit_output_module4[30]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+30]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[30]));
    MUX21X1 U4884(.IN1(head_flit_output_module4[31]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+31]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[31]));
    MUX21X1 U4885(.IN1(head_flit_output_module4[32]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+32]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[32]));
    MUX21X1 U4886(.IN1(head_flit_output_module4[33]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+33]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[33]));
    MUX21X1 U4887(.IN1(head_flit_output_module4[34]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+34]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[34]));
    MUX21X1 U4888(.IN1(head_flit_output_module4[35]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+35]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[35]));
    MUX21X1 U4889(.IN1(head_flit_output_module4[36]), .IN2(int_map_req_v[628:592][in_mod_output_module4[1:0]*37+36]), .S(and2resu1_output_module4) ,.Q(head_flit_output_module4[36]));

    INVX1 U4890 ( .A(head_flit_output_module4[32]), .Y(head_flit_output_module4_32_not_output_module4) );
    AND2X1 U4891 ( .IN1(head_flit_output_module4_32_not_output_module4), .IN2(head_flit_output_module4[33]), .Q(and3resu1_output_module4) );
    NOR4X1 U4892 (.IN1(head_flit_output_module4[29]), .IN2(head_flit_output_module4[28]), .IN3(head_flit_output_module4[27]), .IN4(head_flit_output_module4[26]), .Q(nor23resu1_output_module4) );
    NOR4X1 U4893 (.IN1(head_flit_output_module4[25]), .IN2(head_flit_output_module4[24]), .IN3(head_flit_output_module4[23]), .IN4(head_flit_output_module4[22]), .Q(nor23resu2_output_module4) );
    AND2X1 U4894 ( .IN1(nor23resu1_output_module4), .IN2(nor23resu2_output_module4), .Q(and4resu1_output_module4) );
    NOR2X1 U4895 (.IN1(head_flit_output_module4[33]), .IN2(head_flit_output_module4[32]), .Q(nor23resu3_output_module4) );
    AND2X1 U4896 ( .IN1(nor23resu3_output_module4), .IN2(and4resu1_output_module4), .Q(and5resu1_output_module4) );    
    OR2X1 U4897 (.IN1(and3resu1_output_module4), .IN2(nor23resu3_output_module4), .Q(or12resu12_output_module4) );
    AND2X1 U4898 ( .IN1(ext_resp_v_i[5:4][0]), .IN2(or12resu12_output_module4), .Q(and6resu1_output_module4) );    
    MUX21X1 U4899(.IN1(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]), .IN2(and6resu1_output_module4), .S(and2resu1_output_module4) ,.Q(tail_flit_im_output_module4[vc_channel_output_module4[1:0]]);
    MUX21X1 U4900(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4901(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and2resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    NAND2X1 U4902(.A(_sv2v_jump_output_module4[0]),.B(_sv2v_jump_output_module4[1]),.Y(nand1resu_output_module4));

    AND2X1 U4903 ( .IN1(xor1resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and7resu1) );    
    MUX21X1 U4904(.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4_1[0]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4905(.IN1(_sv2v_jump_output_module4[1]), .IN2(_sv2v_jump_output_module4_1[1]), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    MUX21X1 U4906(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4907(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and7resu1) ,.Q(_sv2v_jump_output_module4[1]);

    HADDX1 U4908 ( .A0(1'b0), .B0(1'b0), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4909 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4910 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4911 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4912 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4913 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4914 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4915 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4916 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4917 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4918 ( .A0(vc_channel_output_module4[0]), .B0(1'b1), .C1(vc_channel_output_module4[1]), .SO(vc_channel_output_module4[0]) );
    HADDX1 U4919 ( .A0(1'b0), .B0(1'b0), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4920 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4921 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );
    HADDX1 U4922 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(in_mod_output_module4[1]), .SO(in_mod_output_module4[0]) );



    BUFX1 U4923(.A(1'b0), .Y(_sv2v_jump_output_module4[0]));
    BUFX1 U4924(.A(1'b0), .Y(_sv2v_jump_output_module4[1]));
    AND2X1 U4925 ( .IN1(xor1resu1_output_module4), .IN2(grant_im_output_module4[i_output_module4[1:0] * 4+:4]), .Q(and8resu1_output_module4) );    
    MUX21X1 U4926(.IN1(vc_ch_act_out_output_module4[0]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[0]);
    MUX21X1 U4927(.IN1(vc_ch_act_out_output_module4[1]), .IN2(i_output_module4[1:0]), .S(and8resu1_output_module4) ,.Q(vc_ch_act_out_output_module4[1]);
    MUX21X1 U4928(.IN1(req_out_output_module4), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(req_out_output_module4);
    MUX21X1 U4929(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4930(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and8resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);
    HADDX1 U4931 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U4932 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    HADDX1 U4933 ( .A0(in_mod_output_module4[0]), .B0(1'b1), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );

    NOR2X1 U4934 (.IN1(_sv2v_jump_output_module4[0]), .IN2(_sv2v_jump_output_module4[1]), .Q(norfinresu1_output_module4) );
    AND2X1 U4935 ( .IN1(norfinresu1_output_module4), .IN2(req_out_output_module4), .Q(and9resu1_output_module4) );    
    HADDX1 U4936 ( .A0(1'b0), .B0(1'b0), .C1(i_output_module4[1]), .SO(i_output_module4[0]) );
    AND2X1 U4937 ( .IN1(and9resu1_output_module4), .IN2(grant_im_output_module4[(vc_ch_act_out_output_module4 * 4) + i_output_module4[1:0]]), .Q(and10resu1_output_module4) );    

    MUX21X1 U4938(.IN1(ext_req_v_o[184:148][3]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+3]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][3]));
    MUX21X1 U4939(.IN1(ext_req_v_o[184:148][4]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+4]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][4]));
    MUX21X1 U4940(.IN1(ext_req_v_o[184:148][5]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+5]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][5]));
    MUX21X1 U4941(.IN1(ext_req_v_o[184:148][6]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+6]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][6]));
    MUX21X1 U4942(.IN1(ext_req_v_o[184:148][7]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+7]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][7]));
    MUX21X1 U4943(.IN1(ext_req_v_o[184:148][8]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+8]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][8]));
    MUX21X1 U4944(.IN1(ext_req_v_o[184:148][9]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+9]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][9]));
    MUX21X1 U4945(.IN1(ext_req_v_o[184:148][10]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+10]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][10]));
    MUX21X1 U4946(.IN1(ext_req_v_o[184:148][11]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+11]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][11]));
    MUX21X1 U4947(.IN1(ext_req_v_o[184:148][12]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+12]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][12]));
    MUX21X1 U4948(.IN1(ext_req_v_o[184:148][13]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+13]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][13]));
    MUX21X1 U4949(.IN1(ext_req_v_o[184:148][14]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+14]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][14]));
    MUX21X1 U4950(.IN1(ext_req_v_o[184:148][15]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+15]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][15]));
    MUX21X1 U4951(.IN1(ext_req_v_o[184:148][16]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+16]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][16]));
    MUX21X1 U4952(.IN1(ext_req_v_o[184:148][17]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+17]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][17]));
    MUX21X1 U4953(.IN1(ext_req_v_o[184:148][18]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+18]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][18]));
    MUX21X1 U4954(.IN1(ext_req_v_o[184:148][19]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+19]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][19]));
    MUX21X1 U4955(.IN1(ext_req_v_o[184:148][20]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+20]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][20]));
    MUX21X1 U4956(.IN1(ext_req_v_o[184:148][21]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+21]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][21]));
    MUX21X1 U4957(.IN1(ext_req_v_o[184:148][22]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+22]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][22]));
    MUX21X1 U4958(.IN1(ext_req_v_o[184:148][23]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+23]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][23]));
    MUX21X1 U4959(.IN1(ext_req_v_o[184:148][24]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+24]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][24]));
    MUX21X1 U4960(.IN1(ext_req_v_o[184:148][25]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+25]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][25]));
    MUX21X1 U4961(.IN1(ext_req_v_o[184:148][26]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+26]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][26]));
    MUX21X1 U4962(.IN1(ext_req_v_o[184:148][27]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+27]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][27]));
    MUX21X1 U4963(.IN1(ext_req_v_o[184:148][28]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+28]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][28]));
    MUX21X1 U4964(.IN1(ext_req_v_o[184:148][29]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+29]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][29]));
    MUX21X1 U4965(.IN1(ext_req_v_o[184:148][30]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+30]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][30]));
    MUX21X1 U4966(.IN1(ext_req_v_o[184:148][31]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+31]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][31]));
    MUX21X1 U4967(.IN1(ext_req_v_o[184:148][32]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+32]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][32]));
    MUX21X1 U4968(.IN1(ext_req_v_o[184:148][33]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+33]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][33]));
    MUX21X1 U4969(.IN1(ext_req_v_o[184:148][34]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+34]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][34]));
    MUX21X1 U4970(.IN1(ext_req_v_o[184:148][35]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+35]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][35]));
    MUX21X1 U4971(.IN1(ext_req_v_o[184:148][36]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37+36]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][36]));

    MUX21X1 U4972(.IN1(ext_req_v_o[184:148][0]), .IN2(int_map_req_v[628:592][i_output_module4[1:0]*37]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][0]);
    MUX21X1 U4973(.IN1(ext_req_v_o[184:148][1]), .IN2(vc_ch_act_out_output_module4[0]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][1]);
    MUX21X1 U4974(.IN1(ext_req_v_o[184:148][2]), .IN2(vc_ch_act_out_output_module4[1]), .S(and10resu1_output_module4) ,.Q(ext_req_v_o[184:148][2]);    
    MUX21X1 U4975(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4976(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b1), .S(and10resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    

    AND2X1 U4977 ( .IN1(and9resu1_output_module4), .IN2(nand1resu_output_module4), .Q(and11resu1_output_module4) );    
    MUX21X1 U4978(.IN1(_sv2v_jump_output_module4[0]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[0]);
    MUX21X1 U4979(.IN1(_sv2v_jump_output_module4[1]), .IN2(1'b0), .S(and11resu1_output_module4) ,.Q(_sv2v_jump_output_module4[1]);    



//router body
	BUFX1 U4980 ( .A(north_recv_req), .Y(ext_req_v_i[0]) );
	BUFX1 U4981 ( .A(north_recv_resp), .Y(ext_resp_v_o[0]) );
	BUFX1 U4982 ( .A(xt_req_v_i[37]), .Y(south_recv_req) );
	BUFX1 U4983 ( .A(south_recv_resp), .Y(ext_resp_v_o[1]) );
	BUFX1 U4984 ( .A(ext_req_v_i[74]), .Y(west_recv_req) );
	BUFX1 U4985 ( .A(west_recv_resp), .Y(ext_resp_v_o[2]) );
	BUFX1 U4986 ( .A(ext_req_v_i[111]), .Y(east_recv_req) );
	BUFX1 U4987 ( .A(east_recv_resp), .Y(ext_resp_v_o[3]) );
	BUFX1 U4988 ( .A(north_send_req), .Y(ext_req_v_o[0]) );
	BUFX1 U4989 ( .A(ext_resp_v_i[0]), .Y(north_send_resp) );
	BUFX1 U4990 ( .A(south_send_req), .Y(ext_req_v_o[37]) );
	BUFX1 U4991 ( .A(ext_resp_v_i[1]), .Y(south_send_resp) );
	BUFX1 U4992 ( .A(west_send_req), .Y(ext_req_v_o[74]) );
	BUFX1 U4993 ( .A(ext_resp_v_i[2]), .Y(west_send_resp) );
	BUFX1 U4994 ( .A(east_send_req), .Y(ext_req_v_o[111]) );
	BUFX1 U4995 ( .A(ext_resp_v_i[3]), .Y(east_send_resp) );
	BUFX1 U4996 ( .A(local_recv_resp), .Y(ext_resp_v_o[4]) );
	BUFX1 U4997 ( .A(ext_req_v_i[148]), .Y(local_recv_req) );
	BUFX1 U4998 ( .A(local_send_req), .Y(ext_req_v_o[148]) );
	BUFX1 U4999 ( .A(ext_resp_v_i[4]), .Y(local_send_resp) );


	MUX21X1 U5000(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[24]) ,.Q(int_map_req_v[0]));
	MUX21X1 U5001(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[24]) ,.Q(int_map_req_v[1]));
	MUX21X1 U5002(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[24]) ,.Q(int_map_req_v[2]));
	MUX21X1 U5003(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[24]) ,.Q(int_map_req_v[3]));
	MUX21X1 U5004(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[24]) ,.Q(int_map_req_v[4]));
	MUX21X1 U5005(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[24]) ,.Q(int_map_req_v[5]));
	MUX21X1 U5006(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[24]) ,.Q(int_map_req_v[6]));
	MUX21X1 U5007(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[24]) ,.Q(int_map_req_v[7]));
	MUX21X1 U5008(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[24]) ,.Q(int_map_req_v[8]));
	MUX21X1 U5009(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[24]) ,.Q(int_map_req_v[9]));
	MUX21X1 U5010(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[24]) ,.Q(int_map_req_v[10]));
	MUX21X1 U5011(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[24]) ,.Q(int_map_req_v[11]));
	MUX21X1 U5012(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[24]) ,.Q(int_map_req_v[12]));
	MUX21X1 U5013(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[24]) ,.Q(int_map_req_v[13]));
	MUX21X1 U5014(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[24]) ,.Q(int_map_req_v[14]));
	MUX21X1 U5015(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[24]) ,.Q(int_map_req_v[15]));
	MUX21X1 U5016(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[24]) ,.Q(int_map_req_v[16]));
	MUX21X1 U5017(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[24]) ,.Q(int_map_req_v[17]));
	MUX21X1 U5018(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[24]) ,.Q(int_map_req_v[18]));
	MUX21X1 U5019(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[24]) ,.Q(int_map_req_v[19]));
	MUX21X1 U5020(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[24]) ,.Q(int_map_req_v[20]));
	MUX21X1 U5021(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[24]) ,.Q(int_map_req_v[21]));
	MUX21X1 U5022(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[24]) ,.Q(int_map_req_v[22]));
	MUX21X1 U5023(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[24]) ,.Q(int_map_req_v[23]));
	MUX21X1 U5024(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[24]) ,.Q(int_map_req_v[24]));
	MUX21X1 U5025(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[24]) ,.Q(int_map_req_v[25]));
	MUX21X1 U5026(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[24]) ,.Q(int_map_req_v[26]));
	MUX21X1 U5027(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[24]) ,.Q(int_map_req_v[27]));
	MUX21X1 U5028(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[24]) ,.Q(int_map_req_v[28]));
	MUX21X1 U5029(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[24]) ,.Q(int_map_req_v[29]));
	MUX21X1 U5030(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[24]) ,.Q(int_map_req_v[30]));
	MUX21X1 U5031(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[24]) ,.Q(int_map_req_v[31]));
	MUX21X1 U5032(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[24]) ,.Q(int_map_req_v[32]));
	MUX21X1 U5033(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[24]) ,.Q(int_map_req_v[33]));
	MUX21X1 U5034(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[24]) ,.Q(int_map_req_v[34]));
	MUX21X1 U5035(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[24]) ,.Q(int_map_req_v[35]));
	MUX21X1 U5036(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[24]) ,.Q(int_map_req_v[36]));
	MUX21X1 U5037(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[19]) ,.Q(int_map_req_v[37]));
	MUX21X1 U5038(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[19]) ,.Q(int_map_req_v[38]));
	MUX21X1 U5039(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[19]) ,.Q(int_map_req_v[39]));
	MUX21X1 U5040(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[19]) ,.Q(int_map_req_v[40]));
	MUX21X1 U5041(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[19]) ,.Q(int_map_req_v[41]));
	MUX21X1 U5042(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[19]) ,.Q(int_map_req_v[42]));
	MUX21X1 U5043(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[19]) ,.Q(int_map_req_v[43]));
	MUX21X1 U5044(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[19]) ,.Q(int_map_req_v[44]));
	MUX21X1 U5045(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[19]) ,.Q(int_map_req_v[45]));
	MUX21X1 U5046(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[19]) ,.Q(int_map_req_v[46]));
	MUX21X1 U5047(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[19]) ,.Q(int_map_req_v[47]));
	MUX21X1 U5048(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[19]) ,.Q(int_map_req_v[48]));
	MUX21X1 U5049(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[19]) ,.Q(int_map_req_v[49]));
	MUX21X1 U5050(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[19]) ,.Q(int_map_req_v[50]));
	MUX21X1 U5051(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[19]) ,.Q(int_map_req_v[51]));
	MUX21X1 U5052(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[19]) ,.Q(int_map_req_v[52]));
	MUX21X1 U5053(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[19]) ,.Q(int_map_req_v[53]));
	MUX21X1 U5054(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[19]) ,.Q(int_map_req_v[54]));
	MUX21X1 U5055(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[19]) ,.Q(int_map_req_v[55]));
	MUX21X1 U5056(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[19]) ,.Q(int_map_req_v[56]));
	MUX21X1 U5057(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[19]) ,.Q(int_map_req_v[57]));
	MUX21X1 U5058(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[19]) ,.Q(int_map_req_v[58]));
	MUX21X1 U5059(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[19]) ,.Q(int_map_req_v[59]));
	MUX21X1 U5060(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[19]) ,.Q(int_map_req_v[60]));
	MUX21X1 U5061(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[19]) ,.Q(int_map_req_v[61]));
	MUX21X1 U5062(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[19]) ,.Q(int_map_req_v[62]));
	MUX21X1 U5063(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[19]) ,.Q(int_map_req_v[63]));
	MUX21X1 U5064(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[19]) ,.Q(int_map_req_v[64]));
	MUX21X1 U5065(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[19]) ,.Q(int_map_req_v[65]));
	MUX21X1 U5066(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[19]) ,.Q(int_map_req_v[66]));
	MUX21X1 U5067(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[19]) ,.Q(int_map_req_v[67]));
	MUX21X1 U5068(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[19]) ,.Q(int_map_req_v[68]));
	MUX21X1 U5069(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[19]) ,.Q(int_map_req_v[69]));
	MUX21X1 U5070(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[19]) ,.Q(int_map_req_v[70]));
	MUX21X1 U5071(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[19]) ,.Q(int_map_req_v[71]));
	MUX21X1 U5072(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[19]) ,.Q(int_map_req_v[72]));
	MUX21X1 U5073(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[19]) ,.Q(int_map_req_v[73]));
	MUX21X1 U5074(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[14]) ,.Q(int_map_req_v[74]));
	MUX21X1 U5075(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[14]) ,.Q(int_map_req_v[75]));
	MUX21X1 U5076(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[14]) ,.Q(int_map_req_v[76]));
	MUX21X1 U5077(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[14]) ,.Q(int_map_req_v[77]));
	MUX21X1 U5078(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[14]) ,.Q(int_map_req_v[78]));
	MUX21X1 U5079(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[14]) ,.Q(int_map_req_v[79]));
	MUX21X1 U5080(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[14]) ,.Q(int_map_req_v[80]));
	MUX21X1 U5081(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[14]) ,.Q(int_map_req_v[81]));
	MUX21X1 U5082(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[14]) ,.Q(int_map_req_v[82]));
	MUX21X1 U5083(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[14]) ,.Q(int_map_req_v[83]));
	MUX21X1 U5084(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[14]) ,.Q(int_map_req_v[84]));
	MUX21X1 U5085(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[14]) ,.Q(int_map_req_v[85]));
	MUX21X1 U5086(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[14]) ,.Q(int_map_req_v[86]));
	MUX21X1 U5087(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[14]) ,.Q(int_map_req_v[87]));
	MUX21X1 U5088(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[14]) ,.Q(int_map_req_v[88]));
	MUX21X1 U5089(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[14]) ,.Q(int_map_req_v[89]));
	MUX21X1 U5090(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[14]) ,.Q(int_map_req_v[90]));
	MUX21X1 U5091(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[14]) ,.Q(int_map_req_v[91]));
	MUX21X1 U5092(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[14]) ,.Q(int_map_req_v[92]));
	MUX21X1 U5093(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[14]) ,.Q(int_map_req_v[93]));
	MUX21X1 U5094(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[14]) ,.Q(int_map_req_v[94]));
	MUX21X1 U5095(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[14]) ,.Q(int_map_req_v[95]));
	MUX21X1 U5096(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[14]) ,.Q(int_map_req_v[96]));
	MUX21X1 U5097(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[14]) ,.Q(int_map_req_v[97]));
	MUX21X1 U5098(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[14]) ,.Q(int_map_req_v[98]));
	MUX21X1 U5099(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[14]) ,.Q(int_map_req_v[99]));
	MUX21X1 U5100(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[14]) ,.Q(int_map_req_v[100]));
	MUX21X1 U5101(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[14]) ,.Q(int_map_req_v[101]));
	MUX21X1 U5102(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[14]) ,.Q(int_map_req_v[102]));
	MUX21X1 U5103(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[14]) ,.Q(int_map_req_v[103]));
	MUX21X1 U5104(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[14]) ,.Q(int_map_req_v[104]));
	MUX21X1 U5105(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[14]) ,.Q(int_map_req_v[105]));
	MUX21X1 U5106(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[14]) ,.Q(int_map_req_v[106]));
	MUX21X1 U5107(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[14]) ,.Q(int_map_req_v[107]));
	MUX21X1 U5108(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[14]) ,.Q(int_map_req_v[108]));
	MUX21X1 U5109(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[14]) ,.Q(int_map_req_v[109]));
	MUX21X1 U5110(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[14]) ,.Q(int_map_req_v[110]));
	MUX21X1 U5111(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[9]) ,.Q(int_map_req_v[111]));
	MUX21X1 U5112(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[9]) ,.Q(int_map_req_v[112]));
	MUX21X1 U5113(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[9]) ,.Q(int_map_req_v[113]));
	MUX21X1 U5114(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[9]) ,.Q(int_map_req_v[114]));
	MUX21X1 U5115(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[9]) ,.Q(int_map_req_v[115]));
	MUX21X1 U5116(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[9]) ,.Q(int_map_req_v[116]));
	MUX21X1 U5117(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[9]) ,.Q(int_map_req_v[117]));
	MUX21X1 U5118(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[9]) ,.Q(int_map_req_v[118]));
	MUX21X1 U5119(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[9]) ,.Q(int_map_req_v[119]));
	MUX21X1 U5120(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[9]) ,.Q(int_map_req_v[120]));
	MUX21X1 U5121(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[9]) ,.Q(int_map_req_v[121]));
	MUX21X1 U5122(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[9]) ,.Q(int_map_req_v[122]));
	MUX21X1 U5123(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[9]) ,.Q(int_map_req_v[123]));
	MUX21X1 U5124(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[9]) ,.Q(int_map_req_v[124]));
	MUX21X1 U5125(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[9]) ,.Q(int_map_req_v[125]));
	MUX21X1 U5126(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[9]) ,.Q(int_map_req_v[126]));
	MUX21X1 U5127(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[9]) ,.Q(int_map_req_v[127]));
	MUX21X1 U5128(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[9]) ,.Q(int_map_req_v[128]));
	MUX21X1 U5129(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[9]) ,.Q(int_map_req_v[129]));
	MUX21X1 U5130(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[9]) ,.Q(int_map_req_v[130]));
	MUX21X1 U5131(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[9]) ,.Q(int_map_req_v[131]));
	MUX21X1 U5132(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[9]) ,.Q(int_map_req_v[132]));
	MUX21X1 U5133(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[9]) ,.Q(int_map_req_v[133]));
	MUX21X1 U5134(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[9]) ,.Q(int_map_req_v[134]));
	MUX21X1 U5135(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[9]) ,.Q(int_map_req_v[135]));
	MUX21X1 U5136(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[9]) ,.Q(int_map_req_v[136]));
	MUX21X1 U5137(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[9]) ,.Q(int_map_req_v[137]));
	MUX21X1 U5138(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[9]) ,.Q(int_map_req_v[138]));
	MUX21X1 U5139(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[9]) ,.Q(int_map_req_v[139]));
	MUX21X1 U5140(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[9]) ,.Q(int_map_req_v[140]));
	MUX21X1 U5141(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[9]) ,.Q(int_map_req_v[141]));
	MUX21X1 U5142(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[9]) ,.Q(int_map_req_v[142]));
	MUX21X1 U5143(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[9]) ,.Q(int_map_req_v[143]));
	MUX21X1 U5144(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[9]) ,.Q(int_map_req_v[144]));
	MUX21X1 U5145(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[9]) ,.Q(int_map_req_v[145]));
	MUX21X1 U5146(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[9]) ,.Q(int_map_req_v[146]));
	MUX21X1 U5147(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[9]) ,.Q(int_map_req_v[147]));
	MUX21X1 U5148(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[3]), .S(int_route_v[9]) ,.Q(int_resp_v[1]));
	MUX21X1 U5149(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[4]), .S(int_route_v[9]) ,.Q(int_resp_v[2]));
	MUX21X1 U5150(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[2]), .S(int_route_v[14]) ,.Q(int_resp_v[2]));
	MUX21X1 U5151(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[3]), .S(int_route_v[14]) ,.Q(int_resp_v[3]));
	MUX21X1 U5152(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[1]), .S(int_route_v[19]) ,.Q(int_resp_v[3]));
	MUX21X1 U5153(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[2]), .S(int_route_v[19]) ,.Q(int_resp_v[4]));
	MUX21X1 U5154(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[0]), .S(int_route_v[24]) ,.Q(int_resp_v[4]));
	MUX21X1 U5155(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[1]), .S(int_route_v[24]) ,.Q(int_resp_v[5]));


	MUX21X1 U5156(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[3]) ,.Q(int_map_req_v[148]));
	MUX21X1 U5157(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[3]) ,.Q(int_map_req_v[149]));
	MUX21X1 U5158(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[3]) ,.Q(int_map_req_v[150]));
	MUX21X1 U5159(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[3]) ,.Q(int_map_req_v[151]));
	MUX21X1 U5160(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[3]) ,.Q(int_map_req_v[152]));
	MUX21X1 U5161(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[3]) ,.Q(int_map_req_v[153]));
	MUX21X1 U5162(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[3]) ,.Q(int_map_req_v[154]));
	MUX21X1 U5163(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[3]) ,.Q(int_map_req_v[155]));
	MUX21X1 U5164(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[3]) ,.Q(int_map_req_v[156]));
	MUX21X1 U5165(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[3]) ,.Q(int_map_req_v[157]));
	MUX21X1 U5166(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[3]) ,.Q(int_map_req_v[158]));
	MUX21X1 U5167(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[3]) ,.Q(int_map_req_v[159]));
	MUX21X1 U5168(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[3]) ,.Q(int_map_req_v[160]));
	MUX21X1 U5169(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[3]) ,.Q(int_map_req_v[161]));
	MUX21X1 U5170(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[3]) ,.Q(int_map_req_v[162]));
	MUX21X1 U5171(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[3]) ,.Q(int_map_req_v[163]));
	MUX21X1 U5172(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[3]) ,.Q(int_map_req_v[164]));
	MUX21X1 U5173(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[3]) ,.Q(int_map_req_v[165]));
	MUX21X1 U5174(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[3]) ,.Q(int_map_req_v[166]));
	MUX21X1 U5175(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[3]) ,.Q(int_map_req_v[167]));
	MUX21X1 U5176(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[3]) ,.Q(int_map_req_v[168]));
	MUX21X1 U5177(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[3]) ,.Q(int_map_req_v[169]));
	MUX21X1 U5178(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[3]) ,.Q(int_map_req_v[170]));
	MUX21X1 U5179(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[3]) ,.Q(int_map_req_v[171]));
	MUX21X1 U5180(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[3]) ,.Q(int_map_req_v[172]));
	MUX21X1 U5181(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[3]) ,.Q(int_map_req_v[173]));
	MUX21X1 U5182(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[3]) ,.Q(int_map_req_v[174]));
	MUX21X1 U5183(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[3]) ,.Q(int_map_req_v[175]));
	MUX21X1 U5184(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[3]) ,.Q(int_map_req_v[176]));
	MUX21X1 U5185(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[3]) ,.Q(int_map_req_v[177]));
	MUX21X1 U5186(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[3]) ,.Q(int_map_req_v[178]));
	MUX21X1 U5187(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[3]) ,.Q(int_map_req_v[179]));
	MUX21X1 U5188(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[3]) ,.Q(int_map_req_v[180]));
	MUX21X1 U5189(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[3]) ,.Q(int_map_req_v[181]));
	MUX21X1 U5190(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[3]) ,.Q(int_map_req_v[182]));
	MUX21X1 U5191(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[3]) ,.Q(int_map_req_v[183]));
	MUX21X1 U5192(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[3]) ,.Q(int_map_req_v[184]));
	MUX21X1 U5193(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[23]) ,.Q(int_map_req_v[185]));
	MUX21X1 U5194(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[23]) ,.Q(int_map_req_v[186]));
	MUX21X1 U5195(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[23]) ,.Q(int_map_req_v[187]));
	MUX21X1 U5196(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[23]) ,.Q(int_map_req_v[188]));
	MUX21X1 U5197(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[23]) ,.Q(int_map_req_v[189]));
	MUX21X1 U5198(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[23]) ,.Q(int_map_req_v[190]));
	MUX21X1 U5199(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[23]) ,.Q(int_map_req_v[191]));
	MUX21X1 U5200(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[23]) ,.Q(int_map_req_v[192]));
	MUX21X1 U5201(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[23]) ,.Q(int_map_req_v[193]));
	MUX21X1 U5202(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[23]) ,.Q(int_map_req_v[194]));
	MUX21X1 U5203(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[23]) ,.Q(int_map_req_v[195]));
	MUX21X1 U5204(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[23]) ,.Q(int_map_req_v[196]));
	MUX21X1 U5205(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[23]) ,.Q(int_map_req_v[197]));
	MUX21X1 U5206(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[23]) ,.Q(int_map_req_v[198]));
	MUX21X1 U5207(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[23]) ,.Q(int_map_req_v[199]));
	MUX21X1 U5208(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[23]) ,.Q(int_map_req_v[200]));
	MUX21X1 U5209(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[23]) ,.Q(int_map_req_v[201]));
	MUX21X1 U5210(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[23]) ,.Q(int_map_req_v[202]));
	MUX21X1 U5211(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[23]) ,.Q(int_map_req_v[203]));
	MUX21X1 U5212(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[23]) ,.Q(int_map_req_v[204]));
	MUX21X1 U5213(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[23]) ,.Q(int_map_req_v[205]));
	MUX21X1 U5214(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[23]) ,.Q(int_map_req_v[206]));
	MUX21X1 U5215(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[23]) ,.Q(int_map_req_v[207]));
	MUX21X1 U5216(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[23]) ,.Q(int_map_req_v[208]));
	MUX21X1 U5217(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[23]) ,.Q(int_map_req_v[209]));
	MUX21X1 U5218(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[23]) ,.Q(int_map_req_v[210]));
	MUX21X1 U5219(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[23]) ,.Q(int_map_req_v[211]));
	MUX21X1 U5220(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[23]) ,.Q(int_map_req_v[212]));
	MUX21X1 U5221(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[23]) ,.Q(int_map_req_v[213]));
	MUX21X1 U5222(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[23]) ,.Q(int_map_req_v[214]));
	MUX21X1 U5223(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[23]) ,.Q(int_map_req_v[215]));
	MUX21X1 U5224(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[23]) ,.Q(int_map_req_v[216]));
	MUX21X1 U5225(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[23]) ,.Q(int_map_req_v[217]));
	MUX21X1 U5226(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[23]) ,.Q(int_map_req_v[218]));
	MUX21X1 U5227(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[23]) ,.Q(int_map_req_v[219]));
	MUX21X1 U5228(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[23]) ,.Q(int_map_req_v[220]));
	MUX21X1 U5229(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[23]) ,.Q(int_map_req_v[221]));
	MUX21X1 U5230(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[18]) ,.Q(int_map_req_v[222]));
	MUX21X1 U5231(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[18]) ,.Q(int_map_req_v[223]));
	MUX21X1 U5232(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[18]) ,.Q(int_map_req_v[224]));
	MUX21X1 U5233(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[18]) ,.Q(int_map_req_v[225]));
	MUX21X1 U5234(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[18]) ,.Q(int_map_req_v[226]));
	MUX21X1 U5235(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[18]) ,.Q(int_map_req_v[227]));
	MUX21X1 U5236(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[18]) ,.Q(int_map_req_v[228]));
	MUX21X1 U5237(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[18]) ,.Q(int_map_req_v[229]));
	MUX21X1 U5238(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[18]) ,.Q(int_map_req_v[230]));
	MUX21X1 U5239(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[18]) ,.Q(int_map_req_v[231]));
	MUX21X1 U5240(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[18]) ,.Q(int_map_req_v[232]));
	MUX21X1 U5241(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[18]) ,.Q(int_map_req_v[233]));
	MUX21X1 U5242(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[18]) ,.Q(int_map_req_v[234]));
	MUX21X1 U5243(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[18]) ,.Q(int_map_req_v[235]));
	MUX21X1 U5244(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[18]) ,.Q(int_map_req_v[236]));
	MUX21X1 U5245(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[18]) ,.Q(int_map_req_v[237]));
	MUX21X1 U5246(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[18]) ,.Q(int_map_req_v[238]));
	MUX21X1 U5247(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[18]) ,.Q(int_map_req_v[239]));
	MUX21X1 U5248(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[18]) ,.Q(int_map_req_v[240]));
	MUX21X1 U5249(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[18]) ,.Q(int_map_req_v[241]));
	MUX21X1 U5250(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[18]) ,.Q(int_map_req_v[242]));
	MUX21X1 U5251(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[18]) ,.Q(int_map_req_v[243]));
	MUX21X1 U5252(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[18]) ,.Q(int_map_req_v[244]));
	MUX21X1 U5253(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[18]) ,.Q(int_map_req_v[245]));
	MUX21X1 U5254(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[18]) ,.Q(int_map_req_v[246]));
	MUX21X1 U5255(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[18]) ,.Q(int_map_req_v[247]));
	MUX21X1 U5256(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[18]) ,.Q(int_map_req_v[248]));
	MUX21X1 U5257(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[18]) ,.Q(int_map_req_v[249]));
	MUX21X1 U5258(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[18]) ,.Q(int_map_req_v[250]));
	MUX21X1 U5259(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[18]) ,.Q(int_map_req_v[251]));
	MUX21X1 U5260(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[18]) ,.Q(int_map_req_v[252]));
	MUX21X1 U5261(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[18]) ,.Q(int_map_req_v[253]));
	MUX21X1 U5262(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[18]) ,.Q(int_map_req_v[254]));
	MUX21X1 U5263(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[18]) ,.Q(int_map_req_v[255]));
	MUX21X1 U5264(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[18]) ,.Q(int_map_req_v[256]));
	MUX21X1 U5265(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[18]) ,.Q(int_map_req_v[257]));
	MUX21X1 U5266(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[18]) ,.Q(int_map_req_v[258]));
	MUX21X1 U5267(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[13]) ,.Q(int_map_req_v[259]));
	MUX21X1 U5268(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[13]) ,.Q(int_map_req_v[260]));
	MUX21X1 U5269(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[13]) ,.Q(int_map_req_v[261]));
	MUX21X1 U5270(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[13]) ,.Q(int_map_req_v[262]));
	MUX21X1 U5271(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[13]) ,.Q(int_map_req_v[263]));
	MUX21X1 U5272(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[13]) ,.Q(int_map_req_v[264]));
	MUX21X1 U5273(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[13]) ,.Q(int_map_req_v[265]));
	MUX21X1 U5274(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[13]) ,.Q(int_map_req_v[266]));
	MUX21X1 U5275(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[13]) ,.Q(int_map_req_v[267]));
	MUX21X1 U5276(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[13]) ,.Q(int_map_req_v[268]));
	MUX21X1 U5277(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[13]) ,.Q(int_map_req_v[269]));
	MUX21X1 U5278(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[13]) ,.Q(int_map_req_v[270]));
	MUX21X1 U5279(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[13]) ,.Q(int_map_req_v[271]));
	MUX21X1 U5280(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[13]) ,.Q(int_map_req_v[272]));
	MUX21X1 U5281(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[13]) ,.Q(int_map_req_v[273]));
	MUX21X1 U5282(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[13]) ,.Q(int_map_req_v[274]));
	MUX21X1 U5283(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[13]) ,.Q(int_map_req_v[275]));
	MUX21X1 U5284(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[13]) ,.Q(int_map_req_v[276]));
	MUX21X1 U5285(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[13]) ,.Q(int_map_req_v[277]));
	MUX21X1 U5286(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[13]) ,.Q(int_map_req_v[278]));
	MUX21X1 U5287(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[13]) ,.Q(int_map_req_v[279]));
	MUX21X1 U5288(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[13]) ,.Q(int_map_req_v[280]));
	MUX21X1 U5289(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[13]) ,.Q(int_map_req_v[281]));
	MUX21X1 U5290(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[13]) ,.Q(int_map_req_v[282]));
	MUX21X1 U5291(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[13]) ,.Q(int_map_req_v[283]));
	MUX21X1 U5292(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[13]) ,.Q(int_map_req_v[284]));
	MUX21X1 U5293(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[13]) ,.Q(int_map_req_v[285]));
	MUX21X1 U5294(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[13]) ,.Q(int_map_req_v[286]));
	MUX21X1 U5295(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[13]) ,.Q(int_map_req_v[287]));
	MUX21X1 U5296(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[13]) ,.Q(int_map_req_v[288]));
	MUX21X1 U5297(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[13]) ,.Q(int_map_req_v[289]));
	MUX21X1 U5298(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[13]) ,.Q(int_map_req_v[290]));
	MUX21X1 U5299(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[13]) ,.Q(int_map_req_v[291]));
	MUX21X1 U5300(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[13]) ,.Q(int_map_req_v[292]));
	MUX21X1 U5301(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[13]) ,.Q(int_map_req_v[293]));
	MUX21X1 U5302(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[13]) ,.Q(int_map_req_v[294]));
	MUX21X1 U5303(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[13]) ,.Q(int_map_req_v[295]));
	MUX21X1 U5304(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[7]), .S(int_route_v[13]) ,.Q(int_resp_v[2]));
	MUX21X1 U5305(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[8]), .S(int_route_v[13]) ,.Q(int_resp_v[3]));
	MUX21X1 U5306(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[6]), .S(int_route_v[18]) ,.Q(int_resp_v[3]));
	MUX21X1 U5307(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[7]), .S(int_route_v[18]) ,.Q(int_resp_v[4]));
	MUX21X1 U5308(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[4]));
	MUX21X1 U5309(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[2]), .S(int_route_v[6]) ,.Q(int_resp_v[5]));
	MUX21X1 U5310(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[0]), .S(int_route_v[4]) ,.Q(int_resp_v[0]));
	MUX21X1 U5311(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));


	MUX21X1 U5312(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[7]) ,.Q(int_map_req_v[296]));
	MUX21X1 U5313(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[7]) ,.Q(int_map_req_v[297]));
	MUX21X1 U5314(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[7]) ,.Q(int_map_req_v[298]));
	MUX21X1 U5315(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[7]) ,.Q(int_map_req_v[299]));
	MUX21X1 U5316(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[7]) ,.Q(int_map_req_v[300]));
	MUX21X1 U5317(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[7]) ,.Q(int_map_req_v[301]));
	MUX21X1 U5318(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[7]) ,.Q(int_map_req_v[302]));
	MUX21X1 U5319(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[7]) ,.Q(int_map_req_v[303]));
	MUX21X1 U5320(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[7]) ,.Q(int_map_req_v[304]));
	MUX21X1 U5321(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[7]) ,.Q(int_map_req_v[305]));
	MUX21X1 U5322(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[7]) ,.Q(int_map_req_v[306]));
	MUX21X1 U5323(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[7]) ,.Q(int_map_req_v[307]));
	MUX21X1 U5324(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[7]) ,.Q(int_map_req_v[308]));
	MUX21X1 U5325(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[7]) ,.Q(int_map_req_v[309]));
	MUX21X1 U5326(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[7]) ,.Q(int_map_req_v[310]));
	MUX21X1 U5327(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[7]) ,.Q(int_map_req_v[311]));
	MUX21X1 U5328(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[7]) ,.Q(int_map_req_v[312]));
	MUX21X1 U5329(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[7]) ,.Q(int_map_req_v[313]));
	MUX21X1 U5330(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[7]) ,.Q(int_map_req_v[314]));
	MUX21X1 U5331(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[7]) ,.Q(int_map_req_v[315]));
	MUX21X1 U5332(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[7]) ,.Q(int_map_req_v[316]));
	MUX21X1 U5333(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[7]) ,.Q(int_map_req_v[317]));
	MUX21X1 U5334(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[7]) ,.Q(int_map_req_v[318]));
	MUX21X1 U5335(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[7]) ,.Q(int_map_req_v[319]));
	MUX21X1 U5336(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[7]) ,.Q(int_map_req_v[320]));
	MUX21X1 U5337(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[7]) ,.Q(int_map_req_v[321]));
	MUX21X1 U5338(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[7]) ,.Q(int_map_req_v[322]));
	MUX21X1 U5339(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[7]) ,.Q(int_map_req_v[323]));
	MUX21X1 U5340(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[7]) ,.Q(int_map_req_v[324]));
	MUX21X1 U5341(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[7]) ,.Q(int_map_req_v[325]));
	MUX21X1 U5342(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[7]) ,.Q(int_map_req_v[326]));
	MUX21X1 U5343(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[7]) ,.Q(int_map_req_v[327]));
	MUX21X1 U5344(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[7]) ,.Q(int_map_req_v[328]));
	MUX21X1 U5345(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[7]) ,.Q(int_map_req_v[329]));
	MUX21X1 U5346(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[7]) ,.Q(int_map_req_v[330]));
	MUX21X1 U5347(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[7]) ,.Q(int_map_req_v[331]));
	MUX21X1 U5348(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[7]) ,.Q(int_map_req_v[332]));
	MUX21X1 U5349(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[2]) ,.Q(int_map_req_v[333]));
	MUX21X1 U5350(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[2]) ,.Q(int_map_req_v[334]));
	MUX21X1 U5351(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[2]) ,.Q(int_map_req_v[335]));
	MUX21X1 U5352(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[2]) ,.Q(int_map_req_v[336]));
	MUX21X1 U5353(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[2]) ,.Q(int_map_req_v[337]));
	MUX21X1 U5354(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[2]) ,.Q(int_map_req_v[338]));
	MUX21X1 U5355(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[2]) ,.Q(int_map_req_v[339]));
	MUX21X1 U5356(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[2]) ,.Q(int_map_req_v[340]));
	MUX21X1 U5357(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[2]) ,.Q(int_map_req_v[341]));
	MUX21X1 U5358(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[2]) ,.Q(int_map_req_v[342]));
	MUX21X1 U5359(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[2]) ,.Q(int_map_req_v[343]));
	MUX21X1 U5360(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[2]) ,.Q(int_map_req_v[344]));
	MUX21X1 U5361(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[2]) ,.Q(int_map_req_v[345]));
	MUX21X1 U5362(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[2]) ,.Q(int_map_req_v[346]));
	MUX21X1 U5363(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[2]) ,.Q(int_map_req_v[347]));
	MUX21X1 U5364(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[2]) ,.Q(int_map_req_v[348]));
	MUX21X1 U5365(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[2]) ,.Q(int_map_req_v[349]));
	MUX21X1 U5366(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[2]) ,.Q(int_map_req_v[350]));
	MUX21X1 U5367(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[2]) ,.Q(int_map_req_v[351]));
	MUX21X1 U5368(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[2]) ,.Q(int_map_req_v[352]));
	MUX21X1 U5369(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[2]) ,.Q(int_map_req_v[353]));
	MUX21X1 U5370(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[2]) ,.Q(int_map_req_v[354]));
	MUX21X1 U5371(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[2]) ,.Q(int_map_req_v[355]));
	MUX21X1 U5372(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[2]) ,.Q(int_map_req_v[356]));
	MUX21X1 U5373(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[2]) ,.Q(int_map_req_v[357]));
	MUX21X1 U5374(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[2]) ,.Q(int_map_req_v[358]));
	MUX21X1 U5375(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[2]) ,.Q(int_map_req_v[359]));
	MUX21X1 U5376(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[2]) ,.Q(int_map_req_v[360]));
	MUX21X1 U5377(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[2]) ,.Q(int_map_req_v[361]));
	MUX21X1 U5378(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[2]) ,.Q(int_map_req_v[362]));
	MUX21X1 U5379(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[2]) ,.Q(int_map_req_v[363]));
	MUX21X1 U5380(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[2]) ,.Q(int_map_req_v[364]));
	MUX21X1 U5381(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[2]) ,.Q(int_map_req_v[365]));
	MUX21X1 U5382(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[2]) ,.Q(int_map_req_v[366]));
	MUX21X1 U5383(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[2]) ,.Q(int_map_req_v[367]));
	MUX21X1 U5384(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[2]) ,.Q(int_map_req_v[368]));
	MUX21X1 U5385(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[2]) ,.Q(int_map_req_v[369]));
	MUX21X1 U5386(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[22]) ,.Q(int_map_req_v[370]));
	MUX21X1 U5387(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[22]) ,.Q(int_map_req_v[371]));
	MUX21X1 U5388(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[22]) ,.Q(int_map_req_v[372]));
	MUX21X1 U5389(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[22]) ,.Q(int_map_req_v[373]));
	MUX21X1 U5390(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[22]) ,.Q(int_map_req_v[374]));
	MUX21X1 U5391(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[22]) ,.Q(int_map_req_v[375]));
	MUX21X1 U5392(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[22]) ,.Q(int_map_req_v[376]));
	MUX21X1 U5393(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[22]) ,.Q(int_map_req_v[377]));
	MUX21X1 U5394(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[22]) ,.Q(int_map_req_v[378]));
	MUX21X1 U5395(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[22]) ,.Q(int_map_req_v[379]));
	MUX21X1 U5396(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[22]) ,.Q(int_map_req_v[380]));
	MUX21X1 U5397(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[22]) ,.Q(int_map_req_v[381]));
	MUX21X1 U5398(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[22]) ,.Q(int_map_req_v[382]));
	MUX21X1 U5399(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[22]) ,.Q(int_map_req_v[383]));
	MUX21X1 U5400(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[22]) ,.Q(int_map_req_v[384]));
	MUX21X1 U5401(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[22]) ,.Q(int_map_req_v[385]));
	MUX21X1 U5402(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[22]) ,.Q(int_map_req_v[386]));
	MUX21X1 U5403(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[22]) ,.Q(int_map_req_v[387]));
	MUX21X1 U5404(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[22]) ,.Q(int_map_req_v[388]));
	MUX21X1 U5405(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[22]) ,.Q(int_map_req_v[389]));
	MUX21X1 U5406(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[22]) ,.Q(int_map_req_v[390]));
	MUX21X1 U5407(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[22]) ,.Q(int_map_req_v[391]));
	MUX21X1 U5408(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[22]) ,.Q(int_map_req_v[392]));
	MUX21X1 U5409(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[22]) ,.Q(int_map_req_v[393]));
	MUX21X1 U5410(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[22]) ,.Q(int_map_req_v[394]));
	MUX21X1 U5411(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[22]) ,.Q(int_map_req_v[395]));
	MUX21X1 U5412(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[22]) ,.Q(int_map_req_v[396]));
	MUX21X1 U5413(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[22]) ,.Q(int_map_req_v[397]));
	MUX21X1 U5414(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[22]) ,.Q(int_map_req_v[398]));
	MUX21X1 U5415(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[22]) ,.Q(int_map_req_v[399]));
	MUX21X1 U5416(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[22]) ,.Q(int_map_req_v[400]));
	MUX21X1 U5417(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[22]) ,.Q(int_map_req_v[401]));
	MUX21X1 U5418(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[22]) ,.Q(int_map_req_v[402]));
	MUX21X1 U5419(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[22]) ,.Q(int_map_req_v[403]));
	MUX21X1 U5420(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[22]) ,.Q(int_map_req_v[404]));
	MUX21X1 U5421(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[22]) ,.Q(int_map_req_v[405]));
	MUX21X1 U5422(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[22]) ,.Q(int_map_req_v[406]));
	MUX21X1 U5423(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[17]) ,.Q(int_map_req_v[407]));
	MUX21X1 U5424(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[17]) ,.Q(int_map_req_v[408]));
	MUX21X1 U5425(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[17]) ,.Q(int_map_req_v[409]));
	MUX21X1 U5426(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[17]) ,.Q(int_map_req_v[410]));
	MUX21X1 U5427(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[17]) ,.Q(int_map_req_v[411]));
	MUX21X1 U5428(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[17]) ,.Q(int_map_req_v[412]));
	MUX21X1 U5429(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[17]) ,.Q(int_map_req_v[413]));
	MUX21X1 U5430(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[17]) ,.Q(int_map_req_v[414]));
	MUX21X1 U5431(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[17]) ,.Q(int_map_req_v[415]));
	MUX21X1 U5432(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[17]) ,.Q(int_map_req_v[416]));
	MUX21X1 U5433(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[17]) ,.Q(int_map_req_v[417]));
	MUX21X1 U5434(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[17]) ,.Q(int_map_req_v[418]));
	MUX21X1 U5435(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[17]) ,.Q(int_map_req_v[419]));
	MUX21X1 U5436(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[17]) ,.Q(int_map_req_v[420]));
	MUX21X1 U5437(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[17]) ,.Q(int_map_req_v[421]));
	MUX21X1 U5438(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[17]) ,.Q(int_map_req_v[422]));
	MUX21X1 U5439(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[17]) ,.Q(int_map_req_v[423]));
	MUX21X1 U5440(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[17]) ,.Q(int_map_req_v[424]));
	MUX21X1 U5441(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[17]) ,.Q(int_map_req_v[425]));
	MUX21X1 U5442(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[17]) ,.Q(int_map_req_v[426]));
	MUX21X1 U5443(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[17]) ,.Q(int_map_req_v[427]));
	MUX21X1 U5444(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[17]) ,.Q(int_map_req_v[428]));
	MUX21X1 U5445(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[17]) ,.Q(int_map_req_v[429]));
	MUX21X1 U5446(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[17]) ,.Q(int_map_req_v[430]));
	MUX21X1 U5447(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[17]) ,.Q(int_map_req_v[431]));
	MUX21X1 U5448(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[17]) ,.Q(int_map_req_v[432]));
	MUX21X1 U5449(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[17]) ,.Q(int_map_req_v[433]));
	MUX21X1 U5450(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[17]) ,.Q(int_map_req_v[434]));
	MUX21X1 U5451(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[17]) ,.Q(int_map_req_v[435]));
	MUX21X1 U5452(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[17]) ,.Q(int_map_req_v[436]));
	MUX21X1 U5453(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[17]) ,.Q(int_map_req_v[437]));
	MUX21X1 U5454(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[17]) ,.Q(int_map_req_v[438]));
	MUX21X1 U5455(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[17]) ,.Q(int_map_req_v[439]));
	MUX21X1 U5456(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[17]) ,.Q(int_map_req_v[440]));
	MUX21X1 U5457(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[17]) ,.Q(int_map_req_v[441]));
	MUX21X1 U5458(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[17]) ,.Q(int_map_req_v[442]));
	MUX21X1 U5459(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[17]) ,.Q(int_map_req_v[443]));
	MUX21X1 U5460(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[11]), .S(int_route_v[17]) ,.Q(int_resp_v[3]));
	MUX21X1 U5461(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[12]), .S(int_route_v[17]) ,.Q(int_resp_v[4]));
	MUX21X1 U5462(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[10]), .S(int_route_v[22]) ,.Q(int_resp_v[4]));
	MUX21X1 U5463(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[11]), .S(int_route_v[22]) ,.Q(int_resp_v[5]));
	MUX21X1 U5464(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[9]), .S(int_route_v[2]) ,.Q(int_resp_v[0]));
	MUX21X1 U5465(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[10]), .S(int_route_v[2]) ,.Q(int_resp_v[1]));
	MUX21X1 U5466(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[8]), .S(int_route_v[7]) ,.Q(int_resp_v[1]));
	MUX21X1 U5467(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[9]), .S(int_route_v[7]) ,.Q(int_resp_v[2]));

	MUX21X1 U5468(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[11]) ,.Q(int_map_req_v[444]));
	MUX21X1 U5469(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[11]) ,.Q(int_map_req_v[445]));
	MUX21X1 U5470(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[11]) ,.Q(int_map_req_v[446]));
	MUX21X1 U5471(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[11]) ,.Q(int_map_req_v[447]));
	MUX21X1 U5472(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[11]) ,.Q(int_map_req_v[448]));
	MUX21X1 U5473(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[11]) ,.Q(int_map_req_v[449]));
	MUX21X1 U5474(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[11]) ,.Q(int_map_req_v[450]));
	MUX21X1 U5475(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[11]) ,.Q(int_map_req_v[451]));
	MUX21X1 U5476(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[11]) ,.Q(int_map_req_v[452]));
	MUX21X1 U5477(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[11]) ,.Q(int_map_req_v[453]));
	MUX21X1 U5478(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[11]) ,.Q(int_map_req_v[454]));
	MUX21X1 U5479(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[11]) ,.Q(int_map_req_v[455]));
	MUX21X1 U5480(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[11]) ,.Q(int_map_req_v[456]));
	MUX21X1 U5481(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[11]) ,.Q(int_map_req_v[457]));
	MUX21X1 U5482(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[11]) ,.Q(int_map_req_v[458]));
	MUX21X1 U5483(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[11]) ,.Q(int_map_req_v[459]));
	MUX21X1 U5484(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[11]) ,.Q(int_map_req_v[460]));
	MUX21X1 U5485(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[11]) ,.Q(int_map_req_v[461]));
	MUX21X1 U5486(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[11]) ,.Q(int_map_req_v[462]));
	MUX21X1 U5487(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[11]) ,.Q(int_map_req_v[463]));
	MUX21X1 U5488(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[11]) ,.Q(int_map_req_v[464]));
	MUX21X1 U5489(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[11]) ,.Q(int_map_req_v[465]));
	MUX21X1 U5490(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[11]) ,.Q(int_map_req_v[466]));
	MUX21X1 U5491(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[11]) ,.Q(int_map_req_v[467]));
	MUX21X1 U5492(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[11]) ,.Q(int_map_req_v[468]));
	MUX21X1 U5493(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[11]) ,.Q(int_map_req_v[469]));
	MUX21X1 U5494(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[11]) ,.Q(int_map_req_v[470]));
	MUX21X1 U5495(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[11]) ,.Q(int_map_req_v[471]));
	MUX21X1 U5496(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[11]) ,.Q(int_map_req_v[472]));
	MUX21X1 U5497(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[11]) ,.Q(int_map_req_v[473]));
	MUX21X1 U5498(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[11]) ,.Q(int_map_req_v[474]));
	MUX21X1 U5499(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[11]) ,.Q(int_map_req_v[475]));
	MUX21X1 U5500(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[11]) ,.Q(int_map_req_v[476]));
	MUX21X1 U5501(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[11]) ,.Q(int_map_req_v[477]));
	MUX21X1 U5502(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[11]) ,.Q(int_map_req_v[478]));
	MUX21X1 U5503(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[11]) ,.Q(int_map_req_v[479]));
	MUX21X1 U5504(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[11]) ,.Q(int_map_req_v[480]));
	MUX21X1 U5505(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[6]) ,.Q(int_map_req_v[481]));
	MUX21X1 U5506(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[6]) ,.Q(int_map_req_v[482]));
	MUX21X1 U5507(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[6]) ,.Q(int_map_req_v[483]));
	MUX21X1 U5508(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[6]) ,.Q(int_map_req_v[484]));
	MUX21X1 U5509(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[6]) ,.Q(int_map_req_v[485]));
	MUX21X1 U5510(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[6]) ,.Q(int_map_req_v[486]));
	MUX21X1 U5511(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[6]) ,.Q(int_map_req_v[487]));
	MUX21X1 U5512(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[6]) ,.Q(int_map_req_v[488]));
	MUX21X1 U5513(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[6]) ,.Q(int_map_req_v[489]));
	MUX21X1 U5514(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[6]) ,.Q(int_map_req_v[490]));
	MUX21X1 U5515(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[6]) ,.Q(int_map_req_v[491]));
	MUX21X1 U5516(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[6]) ,.Q(int_map_req_v[492]));
	MUX21X1 U5517(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[6]) ,.Q(int_map_req_v[493]));
	MUX21X1 U5518(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[6]) ,.Q(int_map_req_v[494]));
	MUX21X1 U5519(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[6]) ,.Q(int_map_req_v[495]));
	MUX21X1 U5520(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[6]) ,.Q(int_map_req_v[496]));
	MUX21X1 U5521(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[6]) ,.Q(int_map_req_v[497]));
	MUX21X1 U5522(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[6]) ,.Q(int_map_req_v[498]));
	MUX21X1 U5523(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[6]) ,.Q(int_map_req_v[499]));
	MUX21X1 U5524(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[6]) ,.Q(int_map_req_v[500]));
	MUX21X1 U5525(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[6]) ,.Q(int_map_req_v[501]));
	MUX21X1 U5526(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[6]) ,.Q(int_map_req_v[502]));
	MUX21X1 U5527(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[6]) ,.Q(int_map_req_v[503]));
	MUX21X1 U5528(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[6]) ,.Q(int_map_req_v[504]));
	MUX21X1 U5529(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[6]) ,.Q(int_map_req_v[505]));
	MUX21X1 U5530(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[6]) ,.Q(int_map_req_v[506]));
	MUX21X1 U5531(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[6]) ,.Q(int_map_req_v[507]));
	MUX21X1 U5532(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[6]) ,.Q(int_map_req_v[508]));
	MUX21X1 U5533(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[6]) ,.Q(int_map_req_v[509]));
	MUX21X1 U5534(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[6]) ,.Q(int_map_req_v[510]));
	MUX21X1 U5535(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[6]) ,.Q(int_map_req_v[511]));
	MUX21X1 U5536(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[6]) ,.Q(int_map_req_v[512]));
	MUX21X1 U5537(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[6]) ,.Q(int_map_req_v[513]));
	MUX21X1 U5538(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[6]) ,.Q(int_map_req_v[514]));
	MUX21X1 U5539(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[6]) ,.Q(int_map_req_v[515]));
	MUX21X1 U5540(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[6]) ,.Q(int_map_req_v[516]));
	MUX21X1 U5541(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[6]) ,.Q(int_map_req_v[517]));
	MUX21X1 U5542(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[1]) ,.Q(int_map_req_v[518]));
	MUX21X1 U5543(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[1]) ,.Q(int_map_req_v[519]));
	MUX21X1 U5544(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[1]) ,.Q(int_map_req_v[520]));
	MUX21X1 U5545(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[1]) ,.Q(int_map_req_v[521]));
	MUX21X1 U5546(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[1]) ,.Q(int_map_req_v[522]));
	MUX21X1 U5547(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[1]) ,.Q(int_map_req_v[523]));
	MUX21X1 U5548(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[1]) ,.Q(int_map_req_v[524]));
	MUX21X1 U5549(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[1]) ,.Q(int_map_req_v[525]));
	MUX21X1 U5550(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[1]) ,.Q(int_map_req_v[526]));
	MUX21X1 U5551(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[1]) ,.Q(int_map_req_v[527]));
	MUX21X1 U5552(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[1]) ,.Q(int_map_req_v[528]));
	MUX21X1 U5553(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[1]) ,.Q(int_map_req_v[529]));
	MUX21X1 U5554(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[1]) ,.Q(int_map_req_v[530]));
	MUX21X1 U5555(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[1]) ,.Q(int_map_req_v[531]));
	MUX21X1 U5556(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[1]) ,.Q(int_map_req_v[532]));
	MUX21X1 U5557(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[1]) ,.Q(int_map_req_v[533]));
	MUX21X1 U5558(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[1]) ,.Q(int_map_req_v[534]));
	MUX21X1 U5559(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[1]) ,.Q(int_map_req_v[535]));
	MUX21X1 U5560(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[1]) ,.Q(int_map_req_v[536]));
	MUX21X1 U5561(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[1]) ,.Q(int_map_req_v[537]));
	MUX21X1 U5562(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[1]) ,.Q(int_map_req_v[538]));
	MUX21X1 U5563(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[1]) ,.Q(int_map_req_v[539]));
	MUX21X1 U5564(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[1]) ,.Q(int_map_req_v[540]));
	MUX21X1 U5565(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[1]) ,.Q(int_map_req_v[541]));
	MUX21X1 U5566(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[1]) ,.Q(int_map_req_v[542]));
	MUX21X1 U5567(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[1]) ,.Q(int_map_req_v[543]));
	MUX21X1 U5568(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[1]) ,.Q(int_map_req_v[544]));
	MUX21X1 U5569(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[1]) ,.Q(int_map_req_v[545]));
	MUX21X1 U5570(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[1]) ,.Q(int_map_req_v[546]));
	MUX21X1 U5571(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[1]) ,.Q(int_map_req_v[547]));
	MUX21X1 U5572(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[1]) ,.Q(int_map_req_v[548]));
	MUX21X1 U5573(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[1]) ,.Q(int_map_req_v[549]));
	MUX21X1 U5574(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[1]) ,.Q(int_map_req_v[550]));
	MUX21X1 U5575(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[1]) ,.Q(int_map_req_v[551]));
	MUX21X1 U5576(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[1]) ,.Q(int_map_req_v[552]));
	MUX21X1 U5577(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[1]) ,.Q(int_map_req_v[553]));
	MUX21X1 U5578(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[1]) ,.Q(int_map_req_v[554]));
	MUX21X1 U5579(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[21]) ,.Q(int_map_req_v[555]));
	MUX21X1 U5580(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[21]) ,.Q(int_map_req_v[556]));
	MUX21X1 U5581(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[21]) ,.Q(int_map_req_v[557]));
	MUX21X1 U5582(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[21]) ,.Q(int_map_req_v[558]));
	MUX21X1 U5583(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[21]) ,.Q(int_map_req_v[559]));
	MUX21X1 U5584(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[21]) ,.Q(int_map_req_v[560]));
	MUX21X1 U5585(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[21]) ,.Q(int_map_req_v[561]));
	MUX21X1 U5586(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[21]) ,.Q(int_map_req_v[562]));
	MUX21X1 U5587(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[21]) ,.Q(int_map_req_v[563]));
	MUX21X1 U5588(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[21]) ,.Q(int_map_req_v[564]));
	MUX21X1 U5589(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[21]) ,.Q(int_map_req_v[565]));
	MUX21X1 U5590(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[21]) ,.Q(int_map_req_v[566]));
	MUX21X1 U5591(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[21]) ,.Q(int_map_req_v[567]));
	MUX21X1 U5592(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[21]) ,.Q(int_map_req_v[568]));
	MUX21X1 U5593(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[21]) ,.Q(int_map_req_v[569]));
	MUX21X1 U5594(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[21]) ,.Q(int_map_req_v[570]));
	MUX21X1 U5595(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[21]) ,.Q(int_map_req_v[571]));
	MUX21X1 U5596(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[21]) ,.Q(int_map_req_v[572]));
	MUX21X1 U5597(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[21]) ,.Q(int_map_req_v[573]));
	MUX21X1 U5598(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[21]) ,.Q(int_map_req_v[574]));
	MUX21X1 U5599(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[21]) ,.Q(int_map_req_v[575]));
	MUX21X1 U5600(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[21]) ,.Q(int_map_req_v[576]));
	MUX21X1 U5601(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[21]) ,.Q(int_map_req_v[577]));
	MUX21X1 U5602(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[21]) ,.Q(int_map_req_v[578]));
	MUX21X1 U5603(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[21]) ,.Q(int_map_req_v[579]));
	MUX21X1 U5604(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[21]) ,.Q(int_map_req_v[580]));
	MUX21X1 U5605(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[21]) ,.Q(int_map_req_v[581]));
	MUX21X1 U5606(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[21]) ,.Q(int_map_req_v[582]));
	MUX21X1 U5607(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[21]) ,.Q(int_map_req_v[583]));
	MUX21X1 U5608(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[21]) ,.Q(int_map_req_v[584]));
	MUX21X1 U5609(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[21]) ,.Q(int_map_req_v[585]));
	MUX21X1 U5610(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[21]) ,.Q(int_map_req_v[586]));
	MUX21X1 U5611(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[21]) ,.Q(int_map_req_v[587]));
	MUX21X1 U5612(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[21]) ,.Q(int_map_req_v[588]));
	MUX21X1 U5613(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[21]) ,.Q(int_map_req_v[589]));
	MUX21X1 U5614(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[21]) ,.Q(int_map_req_v[590]));
	MUX21X1 U5615(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[21]) ,.Q(int_map_req_v[591]));
	MUX21X1 U5616(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[15]), .S(int_route_v[21]) ,.Q(int_resp_v[4]));
	MUX21X1 U5617(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[16]), .S(int_route_v[21]) ,.Q(int_resp_v[5]));
	MUX21X1 U5618(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[14]), .S(int_route_v[1]) ,.Q(int_resp_v[0]));
	MUX21X1 U5619(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[15]), .S(int_route_v[1]) ,.Q(int_resp_v[1]));
	MUX21X1 U5620(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[13]), .S(int_route_v[6]) ,.Q(int_resp_v[1]));
	MUX21X1 U5621(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[14]), .S(int_route_v[6]) ,.Q(int_resp_v[2]));
	MUX21X1 U5622(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[12]), .S(int_route_v[11]) ,.Q(int_resp_v[2]));
	MUX21X1 U5623(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[13]), .S(int_route_v[11]) ,.Q(int_resp_v[3]));



	MUX21X1 U5624(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[15]) ,.Q(int_map_req_v[592]));
	MUX21X1 U5625(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[15]) ,.Q(int_map_req_v[593]));
	MUX21X1 U5626(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[15]) ,.Q(int_map_req_v[594]));
	MUX21X1 U5627(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[15]) ,.Q(int_map_req_v[595]));
	MUX21X1 U5628(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[15]) ,.Q(int_map_req_v[596]));
	MUX21X1 U5629(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[15]) ,.Q(int_map_req_v[597]));
	MUX21X1 U5630(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[15]) ,.Q(int_map_req_v[598]));
	MUX21X1 U5631(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[15]) ,.Q(int_map_req_v[599]));
	MUX21X1 U5632(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[15]) ,.Q(int_map_req_v[600]));
	MUX21X1 U5633(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[15]) ,.Q(int_map_req_v[601]));
	MUX21X1 U5634(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[15]) ,.Q(int_map_req_v[602]));
	MUX21X1 U5635(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[15]) ,.Q(int_map_req_v[603]));
	MUX21X1 U5636(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[15]) ,.Q(int_map_req_v[604]));
	MUX21X1 U5637(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[15]) ,.Q(int_map_req_v[605]));
	MUX21X1 U5638(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[15]) ,.Q(int_map_req_v[606]));
	MUX21X1 U5639(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[15]) ,.Q(int_map_req_v[607]));
	MUX21X1 U5640(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[15]) ,.Q(int_map_req_v[608]));
	MUX21X1 U5641(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[15]) ,.Q(int_map_req_v[609]));
	MUX21X1 U5642(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[15]) ,.Q(int_map_req_v[610]));
	MUX21X1 U5643(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[15]) ,.Q(int_map_req_v[611]));
	MUX21X1 U5644(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[15]) ,.Q(int_map_req_v[612]));
	MUX21X1 U5645(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[15]) ,.Q(int_map_req_v[613]));
	MUX21X1 U5646(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[15]) ,.Q(int_map_req_v[614]));
	MUX21X1 U5647(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[15]) ,.Q(int_map_req_v[615]));
	MUX21X1 U5648(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[15]) ,.Q(int_map_req_v[616]));
	MUX21X1 U5649(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[15]) ,.Q(int_map_req_v[617]));
	MUX21X1 U5650(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[15]) ,.Q(int_map_req_v[618]));
	MUX21X1 U5651(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[15]) ,.Q(int_map_req_v[619]));
	MUX21X1 U5652(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[15]) ,.Q(int_map_req_v[620]));
	MUX21X1 U5653(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[15]) ,.Q(int_map_req_v[621]));
	MUX21X1 U5654(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[15]) ,.Q(int_map_req_v[622]));
	MUX21X1 U5655(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[15]) ,.Q(int_map_req_v[623]));
	MUX21X1 U5656(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[15]) ,.Q(int_map_req_v[624]));
	MUX21X1 U5657(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[15]) ,.Q(int_map_req_v[625]));
	MUX21X1 U5658(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[15]) ,.Q(int_map_req_v[626]));
	MUX21X1 U5659(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[15]) ,.Q(int_map_req_v[627]));
	MUX21X1 U5660(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[15]) ,.Q(int_map_req_v[628]));
	MUX21X1 U5661(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[10]) ,.Q(int_map_req_v[629]));
	MUX21X1 U5662(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[10]) ,.Q(int_map_req_v[630]));
	MUX21X1 U5663(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[10]) ,.Q(int_map_req_v[631]));
	MUX21X1 U5664(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[10]) ,.Q(int_map_req_v[632]));
	MUX21X1 U5665(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[10]) ,.Q(int_map_req_v[633]));
	MUX21X1 U5666(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[10]) ,.Q(int_map_req_v[634]));
	MUX21X1 U5667(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[10]) ,.Q(int_map_req_v[635]));
	MUX21X1 U5668(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[10]) ,.Q(int_map_req_v[636]));
	MUX21X1 U5669(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[10]) ,.Q(int_map_req_v[637]));
	MUX21X1 U5670(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[10]) ,.Q(int_map_req_v[638]));
	MUX21X1 U5671(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[10]) ,.Q(int_map_req_v[639]));
	MUX21X1 U5672(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[10]) ,.Q(int_map_req_v[640]));
	MUX21X1 U5673(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[10]) ,.Q(int_map_req_v[641]));
	MUX21X1 U5674(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[10]) ,.Q(int_map_req_v[642]));
	MUX21X1 U5675(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[10]) ,.Q(int_map_req_v[643]));
	MUX21X1 U5676(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[10]) ,.Q(int_map_req_v[644]));
	MUX21X1 U5677(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[10]) ,.Q(int_map_req_v[645]));
	MUX21X1 U5678(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[10]) ,.Q(int_map_req_v[646]));
	MUX21X1 U5679(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[10]) ,.Q(int_map_req_v[647]));
	MUX21X1 U5680(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[10]) ,.Q(int_map_req_v[648]));
	MUX21X1 U5681(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[10]) ,.Q(int_map_req_v[649]));
	MUX21X1 U5682(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[10]) ,.Q(int_map_req_v[650]));
	MUX21X1 U5683(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[10]) ,.Q(int_map_req_v[651]));
	MUX21X1 U5684(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[10]) ,.Q(int_map_req_v[652]));
	MUX21X1 U5685(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[10]) ,.Q(int_map_req_v[653]));
	MUX21X1 U5686(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[10]) ,.Q(int_map_req_v[654]));
	MUX21X1 U5687(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[10]) ,.Q(int_map_req_v[655]));
	MUX21X1 U5688(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[10]) ,.Q(int_map_req_v[656]));
	MUX21X1 U5689(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[10]) ,.Q(int_map_req_v[657]));
	MUX21X1 U5690(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[10]) ,.Q(int_map_req_v[658]));
	MUX21X1 U5691(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[10]) ,.Q(int_map_req_v[659]));
	MUX21X1 U5692(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[10]) ,.Q(int_map_req_v[660]));
	MUX21X1 U5693(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[10]) ,.Q(int_map_req_v[661]));
	MUX21X1 U5694(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[10]) ,.Q(int_map_req_v[662]));
	MUX21X1 U5695(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[10]) ,.Q(int_map_req_v[663]));
	MUX21X1 U5696(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[10]) ,.Q(int_map_req_v[664]));
	MUX21X1 U5697(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[10]) ,.Q(int_map_req_v[665]));
	MUX21X1 U5698(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[5]) ,.Q(int_map_req_v[666]));
	MUX21X1 U5699(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[5]) ,.Q(int_map_req_v[667]));
	MUX21X1 U5700(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[5]) ,.Q(int_map_req_v[668]));
	MUX21X1 U5701(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[5]) ,.Q(int_map_req_v[669]));
	MUX21X1 U5702(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[5]) ,.Q(int_map_req_v[670]));
	MUX21X1 U5703(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[5]) ,.Q(int_map_req_v[671]));
	MUX21X1 U5704(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[5]) ,.Q(int_map_req_v[672]));
	MUX21X1 U5705(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[5]) ,.Q(int_map_req_v[673]));
	MUX21X1 U5706(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[5]) ,.Q(int_map_req_v[674]));
	MUX21X1 U5707(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[5]) ,.Q(int_map_req_v[675]));
	MUX21X1 U5708(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[5]) ,.Q(int_map_req_v[676]));
	MUX21X1 U5709(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[5]) ,.Q(int_map_req_v[677]));
	MUX21X1 U5710(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[5]) ,.Q(int_map_req_v[678]));
	MUX21X1 U5711(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[5]) ,.Q(int_map_req_v[679]));
	MUX21X1 U5712(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[5]) ,.Q(int_map_req_v[680]));
	MUX21X1 U5713(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[5]) ,.Q(int_map_req_v[681]));
	MUX21X1 U5714(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[5]) ,.Q(int_map_req_v[682]));
	MUX21X1 U5715(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[5]) ,.Q(int_map_req_v[683]));
	MUX21X1 U5716(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[5]) ,.Q(int_map_req_v[684]));
	MUX21X1 U5717(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[5]) ,.Q(int_map_req_v[685]));
	MUX21X1 U5718(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[5]) ,.Q(int_map_req_v[686]));
	MUX21X1 U5719(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[5]) ,.Q(int_map_req_v[687]));
	MUX21X1 U5720(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[5]) ,.Q(int_map_req_v[688]));
	MUX21X1 U5721(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[5]) ,.Q(int_map_req_v[689]));
	MUX21X1 U5722(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[5]) ,.Q(int_map_req_v[690]));
	MUX21X1 U5723(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[5]) ,.Q(int_map_req_v[691]));
	MUX21X1 U5724(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[5]) ,.Q(int_map_req_v[692]));
	MUX21X1 U5725(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[5]) ,.Q(int_map_req_v[693]));
	MUX21X1 U5726(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[5]) ,.Q(int_map_req_v[694]));
	MUX21X1 U5727(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[5]) ,.Q(int_map_req_v[695]));
	MUX21X1 U5728(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[5]) ,.Q(int_map_req_v[696]));
	MUX21X1 U5729(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[5]) ,.Q(int_map_req_v[697]));
	MUX21X1 U5730(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[5]) ,.Q(int_map_req_v[698]));
	MUX21X1 U5731(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[5]) ,.Q(int_map_req_v[699]));
	MUX21X1 U5732(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[5]) ,.Q(int_map_req_v[700]));
	MUX21X1 U5733(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[5]) ,.Q(int_map_req_v[701]));
	MUX21X1 U5734(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[5]) ,.Q(int_map_req_v[702]));
	MUX21X1 U5735(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[0]) ,.Q(int_map_req_v[703]));
	MUX21X1 U5736(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[0]) ,.Q(int_map_req_v[704]));
	MUX21X1 U5737(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[0]) ,.Q(int_map_req_v[705]));
	MUX21X1 U5738(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[0]) ,.Q(int_map_req_v[706]));
	MUX21X1 U5739(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[0]) ,.Q(int_map_req_v[707]));
	MUX21X1 U5740(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[0]) ,.Q(int_map_req_v[708]));
	MUX21X1 U5741(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[0]) ,.Q(int_map_req_v[709]));
	MUX21X1 U5742(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[0]) ,.Q(int_map_req_v[710]));
	MUX21X1 U5743(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[0]) ,.Q(int_map_req_v[711]));
	MUX21X1 U5744(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[0]) ,.Q(int_map_req_v[712]));
	MUX21X1 U5745(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[0]) ,.Q(int_map_req_v[713]));
	MUX21X1 U5746(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[0]) ,.Q(int_map_req_v[714]));
	MUX21X1 U5747(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[0]) ,.Q(int_map_req_v[715]));
	MUX21X1 U5748(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[0]) ,.Q(int_map_req_v[716]));
	MUX21X1 U5749(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[0]) ,.Q(int_map_req_v[717]));
	MUX21X1 U5750(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[0]) ,.Q(int_map_req_v[718]));
	MUX21X1 U5751(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[0]) ,.Q(int_map_req_v[719]));
	MUX21X1 U5752(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[0]) ,.Q(int_map_req_v[720]));
	MUX21X1 U5753(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[0]) ,.Q(int_map_req_v[721]));
	MUX21X1 U5754(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[0]) ,.Q(int_map_req_v[722]));
	MUX21X1 U5755(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[0]) ,.Q(int_map_req_v[723]));
	MUX21X1 U5756(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[0]) ,.Q(int_map_req_v[724]));
	MUX21X1 U5757(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[0]) ,.Q(int_map_req_v[725]));
	MUX21X1 U5758(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[0]) ,.Q(int_map_req_v[726]));
	MUX21X1 U5759(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[0]) ,.Q(int_map_req_v[727]));
	MUX21X1 U5760(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[0]) ,.Q(int_map_req_v[728]));
	MUX21X1 U5761(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[0]) ,.Q(int_map_req_v[729]));
	MUX21X1 U5762(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[0]) ,.Q(int_map_req_v[730]));
	MUX21X1 U5763(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[0]) ,.Q(int_map_req_v[731]));
	MUX21X1 U5764(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[0]) ,.Q(int_map_req_v[732]));
	MUX21X1 U5765(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[0]) ,.Q(int_map_req_v[733]));
	MUX21X1 U5766(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[0]) ,.Q(int_map_req_v[734]));
	MUX21X1 U5767(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[0]) ,.Q(int_map_req_v[735]));
	MUX21X1 U5768(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[0]) ,.Q(int_map_req_v[736]));
	MUX21X1 U5769(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[0]) ,.Q(int_map_req_v[737]));
	MUX21X1 U5770(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[0]) ,.Q(int_map_req_v[738]));
	MUX21X1 U5771(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[0]) ,.Q(int_map_req_v[739]));
	MUX21X1 U5772(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[19]), .S(int_route_v[0]) ,.Q(int_resp_v[0]));
	MUX21X1 U5773(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[20]), .S(int_route_v[0]) ,.Q(int_resp_v[1]));
	MUX21X1 U5774(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[18]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));
	MUX21X1 U5775(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[19]), .S(int_route_v[5]) ,.Q(int_resp_v[2]));
	MUX21X1 U5776(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[17]), .S(int_route_v[10]) ,.Q(int_resp_v[2]));
	MUX21X1 U5777(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[18]), .S(int_route_v[10]) ,.Q(int_resp_v[3]));
	MUX21X1 U5778(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[16]), .S(int_route_v[15]) ,.Q(int_resp_v[3]));
	MUX21X1 U5779(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[17]), .S(int_route_v[15]) ,.Q(int_resp_v[4]));
	
endmodule 