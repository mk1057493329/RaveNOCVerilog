module router_ravenoc (clk,arst,north_send,north_recv,south_send,south_recv,west_send,west_recv,east_send,east_recv,local_send,local_recv);

	input clk;
	input arst;
	input north_send;
	input west_recv;
	input east_send;
	input east_recv;
	input north_recv;
	input south_send;
	input south_recv;
	input west_send;
	input local_send;
	input local_recv;
	
	wire south_recv_resp,south_recv_req,south_send_resp,south_send_req,west_recv_resp,west_recv_req,west_send_resp,west_send_req,north_recv_resp,north_recv_req,north_send_resp,north_send_req,east_recv_resp,east_recv_req,east_send_resp,east_send_req,local_recv_resp,local_recv_req,local_send_resp,local_send_req;
	wire [194:0] int_req_v;
	wire [4:0] int_resp_v;
	wire [24:0] int_route_v;
	wire [739:0] int_map_req_v;
	wire [19:0] int_map_resp_v;
	wire [194:0] ext_req_v_i;
	wire [4:0] ext_resp_v_o;
	wire [194:0] ext_req_v_o;
	wire [4:0] ext_resp_v_i;


//input part
	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[36:0]),
		.fin_resp_o(ext_resp_v_o[1:0]),
		.fout_req_o(int_req_v[36:0]),
		.fout_resp_i(int_resp_v[1:0])
	);
	input_router #(
		.ROUTER_X_ID(0),
		.ROUTER_Y_ID(0)
	) u_input_router(
		.clk(clk),
		.arst(arst),
		.flit_req_i(int_req_v[36:0]),
		.router_port_o(int_route_v[4:0])
	);

	
	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[73:37]),
		.fin_resp_o(ext_resp_v_o[2:1]),
		.fout_req_o(int_req_v[73:37]),
		.fout_resp_i(int_resp_v[2:1])
	);
	input_router #(
		.ROUTER_X_ID(0),
		.ROUTER_Y_ID(0)
	) u_input_router(
		.clk(clk),
		.arst(arst),
		.flit_req_i(int_req_v[73:37]),
		.router_port_o(int_route_v[9:5])
	);


	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[110:74]),
		.fin_resp_o(ext_resp_v_o[3:2]),
		.fout_req_o(int_req_v[110:74]),
		.fout_resp_i(int_resp_v[3:2])
	);
	input_router #(
		.ROUTER_X_ID(0),
		.ROUTER_Y_ID(0)
	) u_input_router(
		.clk(clk),
		.arst(arst),
		.flit_req_i(int_req_v[110:74]),
		.router_port_o(int_route_v[14:10])
	);

	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[147:111]),
		.fin_resp_o(ext_resp_v_o[4:3]),
		.fout_req_o(int_req_v[147:111]),
		.fout_resp_i(int_resp_v[4:3])
	);
	input_router #(
		.ROUTER_X_ID(0),
		.ROUTER_Y_ID(0)
	) u_input_router(
		.clk(clk),
		.arst(arst),
		.flit_req_i(int_req_v[147:111]),
		.router_port_o(int_route_v[19:15])
	);


	
	input_datapath u_input_datapath(
		.clk(clk),
		.arst(arst),
		.fin_req_i(ext_req_v_i[184:148]),
		.fin_resp_o(ext_resp_v_o[5:4]),
		.fout_req_o(int_req_v[184:148]),
		.fout_resp_i(int_resp_v[5:4])
	);
	input_router #(
		.ROUTER_X_ID(0),
		.ROUTER_Y_ID(0)
	) u_input_router(
		.clk(clk),
		.arst(arst),
		.flit_req_i(int_req_v[184:148]),
		.router_port_o(int_route_v[24:20])
	);



//output part	
	output_module u_output_north(
		.clk(clk),
		.arst(arst),
		.fin_req_i(int_map_req_v[36:0]),
		.fin_resp_o(int_map_resp_v[3:0]),
		.fout_req_o(ext_req_v_o[36:0]),
		.fout_resp_i(ext_resp_v_i[1:0])
	);
	output_module u_output_south(
		.clk(clk),
		.arst(arst),
		.fin_req_i(int_map_req_v[184:148]),
		.fin_resp_o(int_map_resp_v[7:4]),
		.fout_req_o(ext_req_v_o[73:37]),
		.fout_resp_i(ext_resp_v_i[2:1])
	);
	output_module u_output_west(
		.clk(clk),
		.arst(arst),
		.fin_req_i(int_map_req_v[332:296]),
		.fin_resp_o(int_map_resp_v[11:8]),
		.fout_req_o(ext_req_v_o[110:74]),
		.fout_resp_i(ext_resp_v_i[3:2])
	);
	output_module u_output_east(
		.clk(clk),
		.arst(arst),
		.fin_req_i(int_map_req_v[480:444]),
		.fin_resp_o(int_map_resp_v[15:12]),
		.fout_req_o(ext_req_v_o[147:111]),
		.fout_resp_i(ext_resp_v_i[4:3])
	);
	output_module u_output_local(
		.clk(clk),
		.arst(arst),
		.fin_req_i(int_map_req_v[628:592]),
		.fin_resp_o(int_map_resp_v[19:16]),
		.fout_req_o(ext_req_v_o[184:148]),
		.fout_resp_i(ext_resp_v_i[5:4])
	);



//router body
	BUFX1 U001 ( .A(north_recv_req), .Y(ext_req_v_i[0]) );
	BUFX1 U002 ( .A(north_recv_resp), .Y(ext_resp_v_o[0]) );
	BUFX1 U003 ( .A(xt_req_v_i[37]), .Y(south_recv_req) );
	BUFX1 U004 ( .A(south_recv_resp), .Y(ext_resp_v_o[1]) );
	BUFX1 U005 ( .A(ext_req_v_i[74]), .Y(west_recv_req) );
	BUFX1 U006 ( .A(west_recv_resp), .Y(ext_resp_v_o[2]) );
	BUFX1 U007 ( .A(ext_req_v_i[111]), .Y(east_recv_req) );
	BUFX1 U008 ( .A(east_recv_resp), .Y(ext_resp_v_o[3]) );
	BUFX1 U009 ( .A(north_send_req), .Y(ext_req_v_o[0]) );
	BUFX1 U010 ( .A(ext_resp_v_i[0]), .Y(north_send_resp) );
	BUFX1 U011 ( .A(south_send_req), .Y(ext_req_v_o[37]) );
	BUFX1 U012 ( .A(ext_resp_v_i[1]), .Y(south_send_resp) );
	BUFX1 U013 ( .A(west_send_req), .Y(ext_req_v_o[74]) );
	BUFX1 U014 ( .A(ext_resp_v_i[2]), .Y(west_send_resp) );
	BUFX1 U015 ( .A(east_send_req), .Y(ext_req_v_o[111]) );
	BUFX1 U016 ( .A(ext_resp_v_i[3]), .Y(east_send_resp) );
	BUFX1 U017 ( .A(local_recv_resp), .Y(ext_resp_v_o[4]) );
	BUFX1 U018 ( .A(ext_req_v_i[148]), .Y(local_recv_req) );
	BUFX1 U019 ( .A(local_send_req), .Y(ext_req_v_o[148]) );
	BUFX1 U020 ( .A(ext_resp_v_i[4]), .Y(local_send_resp) );


	MUX21X1 U0(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[24]) ,.Q(int_map_req_v[0]));
	MUX21X1 U1(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[24]) ,.Q(int_map_req_v[1]));
	MUX21X1 U2(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[24]) ,.Q(int_map_req_v[2]));
	MUX21X1 U3(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[24]) ,.Q(int_map_req_v[3]));
	MUX21X1 U4(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[24]) ,.Q(int_map_req_v[4]));
	MUX21X1 U5(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[24]) ,.Q(int_map_req_v[5]));
	MUX21X1 U6(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[24]) ,.Q(int_map_req_v[6]));
	MUX21X1 U7(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[24]) ,.Q(int_map_req_v[7]));
	MUX21X1 U8(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[24]) ,.Q(int_map_req_v[8]));
	MUX21X1 U9(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[24]) ,.Q(int_map_req_v[9]));
	MUX21X1 U10(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[24]) ,.Q(int_map_req_v[10]));
	MUX21X1 U11(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[24]) ,.Q(int_map_req_v[11]));
	MUX21X1 U12(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[24]) ,.Q(int_map_req_v[12]));
	MUX21X1 U13(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[24]) ,.Q(int_map_req_v[13]));
	MUX21X1 U14(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[24]) ,.Q(int_map_req_v[14]));
	MUX21X1 U15(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[24]) ,.Q(int_map_req_v[15]));
	MUX21X1 U16(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[24]) ,.Q(int_map_req_v[16]));
	MUX21X1 U17(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[24]) ,.Q(int_map_req_v[17]));
	MUX21X1 U18(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[24]) ,.Q(int_map_req_v[18]));
	MUX21X1 U19(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[24]) ,.Q(int_map_req_v[19]));
	MUX21X1 U20(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[24]) ,.Q(int_map_req_v[20]));
	MUX21X1 U21(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[24]) ,.Q(int_map_req_v[21]));
	MUX21X1 U22(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[24]) ,.Q(int_map_req_v[22]));
	MUX21X1 U23(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[24]) ,.Q(int_map_req_v[23]));
	MUX21X1 U24(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[24]) ,.Q(int_map_req_v[24]));
	MUX21X1 U25(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[24]) ,.Q(int_map_req_v[25]));
	MUX21X1 U26(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[24]) ,.Q(int_map_req_v[26]));
	MUX21X1 U27(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[24]) ,.Q(int_map_req_v[27]));
	MUX21X1 U28(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[24]) ,.Q(int_map_req_v[28]));
	MUX21X1 U29(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[24]) ,.Q(int_map_req_v[29]));
	MUX21X1 U30(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[24]) ,.Q(int_map_req_v[30]));
	MUX21X1 U31(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[24]) ,.Q(int_map_req_v[31]));
	MUX21X1 U32(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[24]) ,.Q(int_map_req_v[32]));
	MUX21X1 U33(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[24]) ,.Q(int_map_req_v[33]));
	MUX21X1 U34(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[24]) ,.Q(int_map_req_v[34]));
	MUX21X1 U35(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[24]) ,.Q(int_map_req_v[35]));
	MUX21X1 U36(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[24]) ,.Q(int_map_req_v[36]));
	MUX21X1 U37(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[19]) ,.Q(int_map_req_v[37]));
	MUX21X1 U38(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[19]) ,.Q(int_map_req_v[38]));
	MUX21X1 U39(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[19]) ,.Q(int_map_req_v[39]));
	MUX21X1 U40(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[19]) ,.Q(int_map_req_v[40]));
	MUX21X1 U41(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[19]) ,.Q(int_map_req_v[41]));
	MUX21X1 U42(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[19]) ,.Q(int_map_req_v[42]));
	MUX21X1 U43(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[19]) ,.Q(int_map_req_v[43]));
	MUX21X1 U44(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[19]) ,.Q(int_map_req_v[44]));
	MUX21X1 U45(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[19]) ,.Q(int_map_req_v[45]));
	MUX21X1 U46(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[19]) ,.Q(int_map_req_v[46]));
	MUX21X1 U47(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[19]) ,.Q(int_map_req_v[47]));
	MUX21X1 U48(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[19]) ,.Q(int_map_req_v[48]));
	MUX21X1 U49(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[19]) ,.Q(int_map_req_v[49]));
	MUX21X1 U50(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[19]) ,.Q(int_map_req_v[50]));
	MUX21X1 U51(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[19]) ,.Q(int_map_req_v[51]));
	MUX21X1 U52(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[19]) ,.Q(int_map_req_v[52]));
	MUX21X1 U53(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[19]) ,.Q(int_map_req_v[53]));
	MUX21X1 U54(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[19]) ,.Q(int_map_req_v[54]));
	MUX21X1 U55(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[19]) ,.Q(int_map_req_v[55]));
	MUX21X1 U56(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[19]) ,.Q(int_map_req_v[56]));
	MUX21X1 U57(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[19]) ,.Q(int_map_req_v[57]));
	MUX21X1 U58(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[19]) ,.Q(int_map_req_v[58]));
	MUX21X1 U59(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[19]) ,.Q(int_map_req_v[59]));
	MUX21X1 U60(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[19]) ,.Q(int_map_req_v[60]));
	MUX21X1 U61(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[19]) ,.Q(int_map_req_v[61]));
	MUX21X1 U62(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[19]) ,.Q(int_map_req_v[62]));
	MUX21X1 U63(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[19]) ,.Q(int_map_req_v[63]));
	MUX21X1 U64(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[19]) ,.Q(int_map_req_v[64]));
	MUX21X1 U65(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[19]) ,.Q(int_map_req_v[65]));
	MUX21X1 U66(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[19]) ,.Q(int_map_req_v[66]));
	MUX21X1 U67(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[19]) ,.Q(int_map_req_v[67]));
	MUX21X1 U68(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[19]) ,.Q(int_map_req_v[68]));
	MUX21X1 U69(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[19]) ,.Q(int_map_req_v[69]));
	MUX21X1 U70(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[19]) ,.Q(int_map_req_v[70]));
	MUX21X1 U71(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[19]) ,.Q(int_map_req_v[71]));
	MUX21X1 U72(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[19]) ,.Q(int_map_req_v[72]));
	MUX21X1 U73(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[19]) ,.Q(int_map_req_v[73]));
	MUX21X1 U74(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[14]) ,.Q(int_map_req_v[74]));
	MUX21X1 U75(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[14]) ,.Q(int_map_req_v[75]));
	MUX21X1 U76(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[14]) ,.Q(int_map_req_v[76]));
	MUX21X1 U77(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[14]) ,.Q(int_map_req_v[77]));
	MUX21X1 U78(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[14]) ,.Q(int_map_req_v[78]));
	MUX21X1 U79(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[14]) ,.Q(int_map_req_v[79]));
	MUX21X1 U80(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[14]) ,.Q(int_map_req_v[80]));
	MUX21X1 U81(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[14]) ,.Q(int_map_req_v[81]));
	MUX21X1 U82(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[14]) ,.Q(int_map_req_v[82]));
	MUX21X1 U83(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[14]) ,.Q(int_map_req_v[83]));
	MUX21X1 U84(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[14]) ,.Q(int_map_req_v[84]));
	MUX21X1 U85(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[14]) ,.Q(int_map_req_v[85]));
	MUX21X1 U86(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[14]) ,.Q(int_map_req_v[86]));
	MUX21X1 U87(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[14]) ,.Q(int_map_req_v[87]));
	MUX21X1 U88(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[14]) ,.Q(int_map_req_v[88]));
	MUX21X1 U89(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[14]) ,.Q(int_map_req_v[89]));
	MUX21X1 U90(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[14]) ,.Q(int_map_req_v[90]));
	MUX21X1 U91(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[14]) ,.Q(int_map_req_v[91]));
	MUX21X1 U92(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[14]) ,.Q(int_map_req_v[92]));
	MUX21X1 U93(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[14]) ,.Q(int_map_req_v[93]));
	MUX21X1 U94(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[14]) ,.Q(int_map_req_v[94]));
	MUX21X1 U95(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[14]) ,.Q(int_map_req_v[95]));
	MUX21X1 U96(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[14]) ,.Q(int_map_req_v[96]));
	MUX21X1 U97(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[14]) ,.Q(int_map_req_v[97]));
	MUX21X1 U98(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[14]) ,.Q(int_map_req_v[98]));
	MUX21X1 U99(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[14]) ,.Q(int_map_req_v[99]));
	MUX21X1 U100(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[14]) ,.Q(int_map_req_v[100]));
	MUX21X1 U101(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[14]) ,.Q(int_map_req_v[101]));
	MUX21X1 U102(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[14]) ,.Q(int_map_req_v[102]));
	MUX21X1 U103(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[14]) ,.Q(int_map_req_v[103]));
	MUX21X1 U104(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[14]) ,.Q(int_map_req_v[104]));
	MUX21X1 U105(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[14]) ,.Q(int_map_req_v[105]));
	MUX21X1 U106(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[14]) ,.Q(int_map_req_v[106]));
	MUX21X1 U107(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[14]) ,.Q(int_map_req_v[107]));
	MUX21X1 U108(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[14]) ,.Q(int_map_req_v[108]));
	MUX21X1 U109(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[14]) ,.Q(int_map_req_v[109]));
	MUX21X1 U110(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[14]) ,.Q(int_map_req_v[110]));
	MUX21X1 U111(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[9]) ,.Q(int_map_req_v[111]));
	MUX21X1 U112(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[9]) ,.Q(int_map_req_v[112]));
	MUX21X1 U113(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[9]) ,.Q(int_map_req_v[113]));
	MUX21X1 U114(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[9]) ,.Q(int_map_req_v[114]));
	MUX21X1 U115(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[9]) ,.Q(int_map_req_v[115]));
	MUX21X1 U116(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[9]) ,.Q(int_map_req_v[116]));
	MUX21X1 U117(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[9]) ,.Q(int_map_req_v[117]));
	MUX21X1 U118(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[9]) ,.Q(int_map_req_v[118]));
	MUX21X1 U119(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[9]) ,.Q(int_map_req_v[119]));
	MUX21X1 U120(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[9]) ,.Q(int_map_req_v[120]));
	MUX21X1 U121(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[9]) ,.Q(int_map_req_v[121]));
	MUX21X1 U122(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[9]) ,.Q(int_map_req_v[122]));
	MUX21X1 U123(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[9]) ,.Q(int_map_req_v[123]));
	MUX21X1 U124(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[9]) ,.Q(int_map_req_v[124]));
	MUX21X1 U125(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[9]) ,.Q(int_map_req_v[125]));
	MUX21X1 U126(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[9]) ,.Q(int_map_req_v[126]));
	MUX21X1 U127(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[9]) ,.Q(int_map_req_v[127]));
	MUX21X1 U128(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[9]) ,.Q(int_map_req_v[128]));
	MUX21X1 U129(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[9]) ,.Q(int_map_req_v[129]));
	MUX21X1 U130(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[9]) ,.Q(int_map_req_v[130]));
	MUX21X1 U131(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[9]) ,.Q(int_map_req_v[131]));
	MUX21X1 U132(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[9]) ,.Q(int_map_req_v[132]));
	MUX21X1 U133(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[9]) ,.Q(int_map_req_v[133]));
	MUX21X1 U134(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[9]) ,.Q(int_map_req_v[134]));
	MUX21X1 U135(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[9]) ,.Q(int_map_req_v[135]));
	MUX21X1 U136(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[9]) ,.Q(int_map_req_v[136]));
	MUX21X1 U137(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[9]) ,.Q(int_map_req_v[137]));
	MUX21X1 U138(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[9]) ,.Q(int_map_req_v[138]));
	MUX21X1 U139(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[9]) ,.Q(int_map_req_v[139]));
	MUX21X1 U140(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[9]) ,.Q(int_map_req_v[140]));
	MUX21X1 U141(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[9]) ,.Q(int_map_req_v[141]));
	MUX21X1 U142(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[9]) ,.Q(int_map_req_v[142]));
	MUX21X1 U143(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[9]) ,.Q(int_map_req_v[143]));
	MUX21X1 U144(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[9]) ,.Q(int_map_req_v[144]));
	MUX21X1 U145(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[9]) ,.Q(int_map_req_v[145]));
	MUX21X1 U146(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[9]) ,.Q(int_map_req_v[146]));
	MUX21X1 U147(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[9]) ,.Q(int_map_req_v[147]));
	MUX21X1 U01(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[3]), .S(int_route_v[9]) ,.Q(int_resp_v[1]));
	MUX21X1 U02(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[4]), .S(int_route_v[9]) ,.Q(int_resp_v[2]));
	MUX21X1 U03(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[2]), .S(int_route_v[14]) ,.Q(int_resp_v[2]));
	MUX21X1 U04(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[3]), .S(int_route_v[14]) ,.Q(int_resp_v[3]));
	MUX21X1 U05(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[1]), .S(int_route_v[19]) ,.Q(int_resp_v[3]));
	MUX21X1 U06(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[2]), .S(int_route_v[19]) ,.Q(int_resp_v[4]));
	MUX21X1 U07(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[0]), .S(int_route_v[24]) ,.Q(int_resp_v[4]));
	MUX21X1 U08(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[1]), .S(int_route_v[24]) ,.Q(int_resp_v[5]));


	MUX21X1 U148(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[3]) ,.Q(int_map_req_v[148]));
	MUX21X1 U149(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[3]) ,.Q(int_map_req_v[149]));
	MUX21X1 U150(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[3]) ,.Q(int_map_req_v[150]));
	MUX21X1 U151(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[3]) ,.Q(int_map_req_v[151]));
	MUX21X1 U152(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[3]) ,.Q(int_map_req_v[152]));
	MUX21X1 U153(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[3]) ,.Q(int_map_req_v[153]));
	MUX21X1 U154(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[3]) ,.Q(int_map_req_v[154]));
	MUX21X1 U155(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[3]) ,.Q(int_map_req_v[155]));
	MUX21X1 U156(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[3]) ,.Q(int_map_req_v[156]));
	MUX21X1 U157(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[3]) ,.Q(int_map_req_v[157]));
	MUX21X1 U158(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[3]) ,.Q(int_map_req_v[158]));
	MUX21X1 U159(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[3]) ,.Q(int_map_req_v[159]));
	MUX21X1 U160(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[3]) ,.Q(int_map_req_v[160]));
	MUX21X1 U161(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[3]) ,.Q(int_map_req_v[161]));
	MUX21X1 U162(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[3]) ,.Q(int_map_req_v[162]));
	MUX21X1 U163(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[3]) ,.Q(int_map_req_v[163]));
	MUX21X1 U164(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[3]) ,.Q(int_map_req_v[164]));
	MUX21X1 U165(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[3]) ,.Q(int_map_req_v[165]));
	MUX21X1 U166(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[3]) ,.Q(int_map_req_v[166]));
	MUX21X1 U167(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[3]) ,.Q(int_map_req_v[167]));
	MUX21X1 U168(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[3]) ,.Q(int_map_req_v[168]));
	MUX21X1 U169(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[3]) ,.Q(int_map_req_v[169]));
	MUX21X1 U170(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[3]) ,.Q(int_map_req_v[170]));
	MUX21X1 U171(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[3]) ,.Q(int_map_req_v[171]));
	MUX21X1 U172(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[3]) ,.Q(int_map_req_v[172]));
	MUX21X1 U173(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[3]) ,.Q(int_map_req_v[173]));
	MUX21X1 U174(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[3]) ,.Q(int_map_req_v[174]));
	MUX21X1 U175(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[3]) ,.Q(int_map_req_v[175]));
	MUX21X1 U176(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[3]) ,.Q(int_map_req_v[176]));
	MUX21X1 U177(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[3]) ,.Q(int_map_req_v[177]));
	MUX21X1 U178(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[3]) ,.Q(int_map_req_v[178]));
	MUX21X1 U179(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[3]) ,.Q(int_map_req_v[179]));
	MUX21X1 U180(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[3]) ,.Q(int_map_req_v[180]));
	MUX21X1 U181(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[3]) ,.Q(int_map_req_v[181]));
	MUX21X1 U182(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[3]) ,.Q(int_map_req_v[182]));
	MUX21X1 U183(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[3]) ,.Q(int_map_req_v[183]));
	MUX21X1 U184(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[3]) ,.Q(int_map_req_v[184]));
	MUX21X1 U185(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[23]) ,.Q(int_map_req_v[185]));
	MUX21X1 U186(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[23]) ,.Q(int_map_req_v[186]));
	MUX21X1 U187(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[23]) ,.Q(int_map_req_v[187]));
	MUX21X1 U188(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[23]) ,.Q(int_map_req_v[188]));
	MUX21X1 U189(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[23]) ,.Q(int_map_req_v[189]));
	MUX21X1 U190(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[23]) ,.Q(int_map_req_v[190]));
	MUX21X1 U191(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[23]) ,.Q(int_map_req_v[191]));
	MUX21X1 U192(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[23]) ,.Q(int_map_req_v[192]));
	MUX21X1 U193(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[23]) ,.Q(int_map_req_v[193]));
	MUX21X1 U194(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[23]) ,.Q(int_map_req_v[194]));
	MUX21X1 U195(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[23]) ,.Q(int_map_req_v[195]));
	MUX21X1 U196(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[23]) ,.Q(int_map_req_v[196]));
	MUX21X1 U197(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[23]) ,.Q(int_map_req_v[197]));
	MUX21X1 U198(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[23]) ,.Q(int_map_req_v[198]));
	MUX21X1 U199(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[23]) ,.Q(int_map_req_v[199]));
	MUX21X1 U200(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[23]) ,.Q(int_map_req_v[200]));
	MUX21X1 U201(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[23]) ,.Q(int_map_req_v[201]));
	MUX21X1 U202(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[23]) ,.Q(int_map_req_v[202]));
	MUX21X1 U203(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[23]) ,.Q(int_map_req_v[203]));
	MUX21X1 U204(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[23]) ,.Q(int_map_req_v[204]));
	MUX21X1 U205(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[23]) ,.Q(int_map_req_v[205]));
	MUX21X1 U206(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[23]) ,.Q(int_map_req_v[206]));
	MUX21X1 U207(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[23]) ,.Q(int_map_req_v[207]));
	MUX21X1 U208(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[23]) ,.Q(int_map_req_v[208]));
	MUX21X1 U209(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[23]) ,.Q(int_map_req_v[209]));
	MUX21X1 U210(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[23]) ,.Q(int_map_req_v[210]));
	MUX21X1 U211(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[23]) ,.Q(int_map_req_v[211]));
	MUX21X1 U212(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[23]) ,.Q(int_map_req_v[212]));
	MUX21X1 U213(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[23]) ,.Q(int_map_req_v[213]));
	MUX21X1 U214(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[23]) ,.Q(int_map_req_v[214]));
	MUX21X1 U215(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[23]) ,.Q(int_map_req_v[215]));
	MUX21X1 U216(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[23]) ,.Q(int_map_req_v[216]));
	MUX21X1 U217(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[23]) ,.Q(int_map_req_v[217]));
	MUX21X1 U218(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[23]) ,.Q(int_map_req_v[218]));
	MUX21X1 U219(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[23]) ,.Q(int_map_req_v[219]));
	MUX21X1 U220(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[23]) ,.Q(int_map_req_v[220]));
	MUX21X1 U221(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[23]) ,.Q(int_map_req_v[221]));
	MUX21X1 U222(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[18]) ,.Q(int_map_req_v[222]));
	MUX21X1 U223(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[18]) ,.Q(int_map_req_v[223]));
	MUX21X1 U224(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[18]) ,.Q(int_map_req_v[224]));
	MUX21X1 U225(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[18]) ,.Q(int_map_req_v[225]));
	MUX21X1 U226(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[18]) ,.Q(int_map_req_v[226]));
	MUX21X1 U227(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[18]) ,.Q(int_map_req_v[227]));
	MUX21X1 U228(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[18]) ,.Q(int_map_req_v[228]));
	MUX21X1 U229(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[18]) ,.Q(int_map_req_v[229]));
	MUX21X1 U230(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[18]) ,.Q(int_map_req_v[230]));
	MUX21X1 U231(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[18]) ,.Q(int_map_req_v[231]));
	MUX21X1 U232(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[18]) ,.Q(int_map_req_v[232]));
	MUX21X1 U233(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[18]) ,.Q(int_map_req_v[233]));
	MUX21X1 U234(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[18]) ,.Q(int_map_req_v[234]));
	MUX21X1 U235(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[18]) ,.Q(int_map_req_v[235]));
	MUX21X1 U236(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[18]) ,.Q(int_map_req_v[236]));
	MUX21X1 U237(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[18]) ,.Q(int_map_req_v[237]));
	MUX21X1 U238(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[18]) ,.Q(int_map_req_v[238]));
	MUX21X1 U239(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[18]) ,.Q(int_map_req_v[239]));
	MUX21X1 U240(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[18]) ,.Q(int_map_req_v[240]));
	MUX21X1 U241(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[18]) ,.Q(int_map_req_v[241]));
	MUX21X1 U242(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[18]) ,.Q(int_map_req_v[242]));
	MUX21X1 U243(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[18]) ,.Q(int_map_req_v[243]));
	MUX21X1 U244(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[18]) ,.Q(int_map_req_v[244]));
	MUX21X1 U245(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[18]) ,.Q(int_map_req_v[245]));
	MUX21X1 U246(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[18]) ,.Q(int_map_req_v[246]));
	MUX21X1 U247(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[18]) ,.Q(int_map_req_v[247]));
	MUX21X1 U248(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[18]) ,.Q(int_map_req_v[248]));
	MUX21X1 U249(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[18]) ,.Q(int_map_req_v[249]));
	MUX21X1 U250(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[18]) ,.Q(int_map_req_v[250]));
	MUX21X1 U251(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[18]) ,.Q(int_map_req_v[251]));
	MUX21X1 U252(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[18]) ,.Q(int_map_req_v[252]));
	MUX21X1 U253(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[18]) ,.Q(int_map_req_v[253]));
	MUX21X1 U254(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[18]) ,.Q(int_map_req_v[254]));
	MUX21X1 U255(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[18]) ,.Q(int_map_req_v[255]));
	MUX21X1 U256(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[18]) ,.Q(int_map_req_v[256]));
	MUX21X1 U257(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[18]) ,.Q(int_map_req_v[257]));
	MUX21X1 U258(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[18]) ,.Q(int_map_req_v[258]));
	MUX21X1 U259(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[13]) ,.Q(int_map_req_v[259]));
	MUX21X1 U260(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[13]) ,.Q(int_map_req_v[260]));
	MUX21X1 U261(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[13]) ,.Q(int_map_req_v[261]));
	MUX21X1 U262(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[13]) ,.Q(int_map_req_v[262]));
	MUX21X1 U263(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[13]) ,.Q(int_map_req_v[263]));
	MUX21X1 U264(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[13]) ,.Q(int_map_req_v[264]));
	MUX21X1 U265(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[13]) ,.Q(int_map_req_v[265]));
	MUX21X1 U266(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[13]) ,.Q(int_map_req_v[266]));
	MUX21X1 U267(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[13]) ,.Q(int_map_req_v[267]));
	MUX21X1 U268(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[13]) ,.Q(int_map_req_v[268]));
	MUX21X1 U269(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[13]) ,.Q(int_map_req_v[269]));
	MUX21X1 U270(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[13]) ,.Q(int_map_req_v[270]));
	MUX21X1 U271(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[13]) ,.Q(int_map_req_v[271]));
	MUX21X1 U272(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[13]) ,.Q(int_map_req_v[272]));
	MUX21X1 U273(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[13]) ,.Q(int_map_req_v[273]));
	MUX21X1 U274(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[13]) ,.Q(int_map_req_v[274]));
	MUX21X1 U275(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[13]) ,.Q(int_map_req_v[275]));
	MUX21X1 U276(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[13]) ,.Q(int_map_req_v[276]));
	MUX21X1 U277(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[13]) ,.Q(int_map_req_v[277]));
	MUX21X1 U278(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[13]) ,.Q(int_map_req_v[278]));
	MUX21X1 U279(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[13]) ,.Q(int_map_req_v[279]));
	MUX21X1 U280(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[13]) ,.Q(int_map_req_v[280]));
	MUX21X1 U281(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[13]) ,.Q(int_map_req_v[281]));
	MUX21X1 U282(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[13]) ,.Q(int_map_req_v[282]));
	MUX21X1 U283(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[13]) ,.Q(int_map_req_v[283]));
	MUX21X1 U284(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[13]) ,.Q(int_map_req_v[284]));
	MUX21X1 U285(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[13]) ,.Q(int_map_req_v[285]));
	MUX21X1 U286(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[13]) ,.Q(int_map_req_v[286]));
	MUX21X1 U287(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[13]) ,.Q(int_map_req_v[287]));
	MUX21X1 U288(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[13]) ,.Q(int_map_req_v[288]));
	MUX21X1 U289(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[13]) ,.Q(int_map_req_v[289]));
	MUX21X1 U290(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[13]) ,.Q(int_map_req_v[290]));
	MUX21X1 U291(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[13]) ,.Q(int_map_req_v[291]));
	MUX21X1 U292(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[13]) ,.Q(int_map_req_v[292]));
	MUX21X1 U293(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[13]) ,.Q(int_map_req_v[293]));
	MUX21X1 U294(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[13]) ,.Q(int_map_req_v[294]));
	MUX21X1 U295(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[13]) ,.Q(int_map_req_v[295]));
	MUX21X1 U09(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[7]), .S(int_route_v[13]) ,.Q(int_resp_v[2]));
	MUX21X1 U10(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[8]), .S(int_route_v[13]) ,.Q(int_resp_v[3]));
	MUX21X1 U11(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[6]), .S(int_route_v[18]) ,.Q(int_resp_v[3]));
	MUX21X1 U12(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[7]), .S(int_route_v[18]) ,.Q(int_resp_v[4]));
	MUX21X1 U13(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[4]));
	MUX21X1 U14(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[2]), .S(int_route_v[6]) ,.Q(int_resp_v[5]));
	MUX21X1 U15(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[0]), .S(int_route_v[4]) ,.Q(int_resp_v[0]));
	MUX21X1 U16(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[1]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));


	MUX21X1 U296(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[7]) ,.Q(int_map_req_v[296]));
	MUX21X1 U297(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[7]) ,.Q(int_map_req_v[297]));
	MUX21X1 U298(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[7]) ,.Q(int_map_req_v[298]));
	MUX21X1 U299(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[7]) ,.Q(int_map_req_v[299]));
	MUX21X1 U300(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[7]) ,.Q(int_map_req_v[300]));
	MUX21X1 U301(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[7]) ,.Q(int_map_req_v[301]));
	MUX21X1 U302(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[7]) ,.Q(int_map_req_v[302]));
	MUX21X1 U303(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[7]) ,.Q(int_map_req_v[303]));
	MUX21X1 U304(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[7]) ,.Q(int_map_req_v[304]));
	MUX21X1 U305(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[7]) ,.Q(int_map_req_v[305]));
	MUX21X1 U306(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[7]) ,.Q(int_map_req_v[306]));
	MUX21X1 U307(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[7]) ,.Q(int_map_req_v[307]));
	MUX21X1 U308(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[7]) ,.Q(int_map_req_v[308]));
	MUX21X1 U309(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[7]) ,.Q(int_map_req_v[309]));
	MUX21X1 U310(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[7]) ,.Q(int_map_req_v[310]));
	MUX21X1 U311(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[7]) ,.Q(int_map_req_v[311]));
	MUX21X1 U312(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[7]) ,.Q(int_map_req_v[312]));
	MUX21X1 U313(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[7]) ,.Q(int_map_req_v[313]));
	MUX21X1 U314(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[7]) ,.Q(int_map_req_v[314]));
	MUX21X1 U315(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[7]) ,.Q(int_map_req_v[315]));
	MUX21X1 U316(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[7]) ,.Q(int_map_req_v[316]));
	MUX21X1 U317(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[7]) ,.Q(int_map_req_v[317]));
	MUX21X1 U318(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[7]) ,.Q(int_map_req_v[318]));
	MUX21X1 U319(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[7]) ,.Q(int_map_req_v[319]));
	MUX21X1 U320(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[7]) ,.Q(int_map_req_v[320]));
	MUX21X1 U321(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[7]) ,.Q(int_map_req_v[321]));
	MUX21X1 U322(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[7]) ,.Q(int_map_req_v[322]));
	MUX21X1 U323(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[7]) ,.Q(int_map_req_v[323]));
	MUX21X1 U324(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[7]) ,.Q(int_map_req_v[324]));
	MUX21X1 U325(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[7]) ,.Q(int_map_req_v[325]));
	MUX21X1 U326(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[7]) ,.Q(int_map_req_v[326]));
	MUX21X1 U327(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[7]) ,.Q(int_map_req_v[327]));
	MUX21X1 U328(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[7]) ,.Q(int_map_req_v[328]));
	MUX21X1 U329(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[7]) ,.Q(int_map_req_v[329]));
	MUX21X1 U330(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[7]) ,.Q(int_map_req_v[330]));
	MUX21X1 U331(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[7]) ,.Q(int_map_req_v[331]));
	MUX21X1 U332(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[7]) ,.Q(int_map_req_v[332]));
	MUX21X1 U333(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[2]) ,.Q(int_map_req_v[333]));
	MUX21X1 U334(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[2]) ,.Q(int_map_req_v[334]));
	MUX21X1 U335(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[2]) ,.Q(int_map_req_v[335]));
	MUX21X1 U336(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[2]) ,.Q(int_map_req_v[336]));
	MUX21X1 U337(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[2]) ,.Q(int_map_req_v[337]));
	MUX21X1 U338(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[2]) ,.Q(int_map_req_v[338]));
	MUX21X1 U339(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[2]) ,.Q(int_map_req_v[339]));
	MUX21X1 U340(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[2]) ,.Q(int_map_req_v[340]));
	MUX21X1 U341(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[2]) ,.Q(int_map_req_v[341]));
	MUX21X1 U342(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[2]) ,.Q(int_map_req_v[342]));
	MUX21X1 U343(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[2]) ,.Q(int_map_req_v[343]));
	MUX21X1 U344(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[2]) ,.Q(int_map_req_v[344]));
	MUX21X1 U345(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[2]) ,.Q(int_map_req_v[345]));
	MUX21X1 U346(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[2]) ,.Q(int_map_req_v[346]));
	MUX21X1 U347(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[2]) ,.Q(int_map_req_v[347]));
	MUX21X1 U348(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[2]) ,.Q(int_map_req_v[348]));
	MUX21X1 U349(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[2]) ,.Q(int_map_req_v[349]));
	MUX21X1 U350(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[2]) ,.Q(int_map_req_v[350]));
	MUX21X1 U351(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[2]) ,.Q(int_map_req_v[351]));
	MUX21X1 U352(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[2]) ,.Q(int_map_req_v[352]));
	MUX21X1 U353(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[2]) ,.Q(int_map_req_v[353]));
	MUX21X1 U354(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[2]) ,.Q(int_map_req_v[354]));
	MUX21X1 U355(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[2]) ,.Q(int_map_req_v[355]));
	MUX21X1 U356(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[2]) ,.Q(int_map_req_v[356]));
	MUX21X1 U357(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[2]) ,.Q(int_map_req_v[357]));
	MUX21X1 U358(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[2]) ,.Q(int_map_req_v[358]));
	MUX21X1 U359(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[2]) ,.Q(int_map_req_v[359]));
	MUX21X1 U360(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[2]) ,.Q(int_map_req_v[360]));
	MUX21X1 U361(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[2]) ,.Q(int_map_req_v[361]));
	MUX21X1 U362(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[2]) ,.Q(int_map_req_v[362]));
	MUX21X1 U363(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[2]) ,.Q(int_map_req_v[363]));
	MUX21X1 U364(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[2]) ,.Q(int_map_req_v[364]));
	MUX21X1 U365(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[2]) ,.Q(int_map_req_v[365]));
	MUX21X1 U366(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[2]) ,.Q(int_map_req_v[366]));
	MUX21X1 U367(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[2]) ,.Q(int_map_req_v[367]));
	MUX21X1 U368(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[2]) ,.Q(int_map_req_v[368]));
	MUX21X1 U369(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[2]) ,.Q(int_map_req_v[369]));
	MUX21X1 U370(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[22]) ,.Q(int_map_req_v[370]));
	MUX21X1 U371(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[22]) ,.Q(int_map_req_v[371]));
	MUX21X1 U372(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[22]) ,.Q(int_map_req_v[372]));
	MUX21X1 U373(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[22]) ,.Q(int_map_req_v[373]));
	MUX21X1 U374(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[22]) ,.Q(int_map_req_v[374]));
	MUX21X1 U375(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[22]) ,.Q(int_map_req_v[375]));
	MUX21X1 U376(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[22]) ,.Q(int_map_req_v[376]));
	MUX21X1 U377(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[22]) ,.Q(int_map_req_v[377]));
	MUX21X1 U378(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[22]) ,.Q(int_map_req_v[378]));
	MUX21X1 U379(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[22]) ,.Q(int_map_req_v[379]));
	MUX21X1 U380(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[22]) ,.Q(int_map_req_v[380]));
	MUX21X1 U381(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[22]) ,.Q(int_map_req_v[381]));
	MUX21X1 U382(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[22]) ,.Q(int_map_req_v[382]));
	MUX21X1 U383(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[22]) ,.Q(int_map_req_v[383]));
	MUX21X1 U384(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[22]) ,.Q(int_map_req_v[384]));
	MUX21X1 U385(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[22]) ,.Q(int_map_req_v[385]));
	MUX21X1 U386(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[22]) ,.Q(int_map_req_v[386]));
	MUX21X1 U387(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[22]) ,.Q(int_map_req_v[387]));
	MUX21X1 U388(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[22]) ,.Q(int_map_req_v[388]));
	MUX21X1 U389(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[22]) ,.Q(int_map_req_v[389]));
	MUX21X1 U390(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[22]) ,.Q(int_map_req_v[390]));
	MUX21X1 U391(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[22]) ,.Q(int_map_req_v[391]));
	MUX21X1 U392(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[22]) ,.Q(int_map_req_v[392]));
	MUX21X1 U393(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[22]) ,.Q(int_map_req_v[393]));
	MUX21X1 U394(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[22]) ,.Q(int_map_req_v[394]));
	MUX21X1 U395(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[22]) ,.Q(int_map_req_v[395]));
	MUX21X1 U396(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[22]) ,.Q(int_map_req_v[396]));
	MUX21X1 U397(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[22]) ,.Q(int_map_req_v[397]));
	MUX21X1 U398(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[22]) ,.Q(int_map_req_v[398]));
	MUX21X1 U399(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[22]) ,.Q(int_map_req_v[399]));
	MUX21X1 U400(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[22]) ,.Q(int_map_req_v[400]));
	MUX21X1 U401(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[22]) ,.Q(int_map_req_v[401]));
	MUX21X1 U402(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[22]) ,.Q(int_map_req_v[402]));
	MUX21X1 U403(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[22]) ,.Q(int_map_req_v[403]));
	MUX21X1 U404(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[22]) ,.Q(int_map_req_v[404]));
	MUX21X1 U405(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[22]) ,.Q(int_map_req_v[405]));
	MUX21X1 U406(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[22]) ,.Q(int_map_req_v[406]));
	MUX21X1 U407(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[17]) ,.Q(int_map_req_v[407]));
	MUX21X1 U408(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[17]) ,.Q(int_map_req_v[408]));
	MUX21X1 U409(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[17]) ,.Q(int_map_req_v[409]));
	MUX21X1 U410(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[17]) ,.Q(int_map_req_v[410]));
	MUX21X1 U411(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[17]) ,.Q(int_map_req_v[411]));
	MUX21X1 U412(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[17]) ,.Q(int_map_req_v[412]));
	MUX21X1 U413(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[17]) ,.Q(int_map_req_v[413]));
	MUX21X1 U414(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[17]) ,.Q(int_map_req_v[414]));
	MUX21X1 U415(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[17]) ,.Q(int_map_req_v[415]));
	MUX21X1 U416(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[17]) ,.Q(int_map_req_v[416]));
	MUX21X1 U417(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[17]) ,.Q(int_map_req_v[417]));
	MUX21X1 U418(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[17]) ,.Q(int_map_req_v[418]));
	MUX21X1 U419(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[17]) ,.Q(int_map_req_v[419]));
	MUX21X1 U420(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[17]) ,.Q(int_map_req_v[420]));
	MUX21X1 U421(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[17]) ,.Q(int_map_req_v[421]));
	MUX21X1 U422(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[17]) ,.Q(int_map_req_v[422]));
	MUX21X1 U423(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[17]) ,.Q(int_map_req_v[423]));
	MUX21X1 U424(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[17]) ,.Q(int_map_req_v[424]));
	MUX21X1 U425(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[17]) ,.Q(int_map_req_v[425]));
	MUX21X1 U426(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[17]) ,.Q(int_map_req_v[426]));
	MUX21X1 U427(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[17]) ,.Q(int_map_req_v[427]));
	MUX21X1 U428(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[17]) ,.Q(int_map_req_v[428]));
	MUX21X1 U429(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[17]) ,.Q(int_map_req_v[429]));
	MUX21X1 U430(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[17]) ,.Q(int_map_req_v[430]));
	MUX21X1 U431(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[17]) ,.Q(int_map_req_v[431]));
	MUX21X1 U432(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[17]) ,.Q(int_map_req_v[432]));
	MUX21X1 U433(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[17]) ,.Q(int_map_req_v[433]));
	MUX21X1 U434(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[17]) ,.Q(int_map_req_v[434]));
	MUX21X1 U435(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[17]) ,.Q(int_map_req_v[435]));
	MUX21X1 U436(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[17]) ,.Q(int_map_req_v[436]));
	MUX21X1 U437(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[17]) ,.Q(int_map_req_v[437]));
	MUX21X1 U438(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[17]) ,.Q(int_map_req_v[438]));
	MUX21X1 U439(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[17]) ,.Q(int_map_req_v[439]));
	MUX21X1 U440(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[17]) ,.Q(int_map_req_v[440]));
	MUX21X1 U441(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[17]) ,.Q(int_map_req_v[441]));
	MUX21X1 U442(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[17]) ,.Q(int_map_req_v[442]));
	MUX21X1 U443(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[17]) ,.Q(int_map_req_v[443]));
	MUX21X1 U17(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[11]), .S(int_route_v[17]) ,.Q(int_resp_v[3]));
	MUX21X1 U18(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[12]), .S(int_route_v[17]) ,.Q(int_resp_v[4]));
	MUX21X1 U19(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[10]), .S(int_route_v[22]) ,.Q(int_resp_v[4]));
	MUX21X1 U20(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[11]), .S(int_route_v[22]) ,.Q(int_resp_v[5]));
	MUX21X1 U21(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[9]), .S(int_route_v[2]) ,.Q(int_resp_v[0]));
	MUX21X1 U22(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[10]), .S(int_route_v[2]) ,.Q(int_resp_v[1]));
	MUX21X1 U23(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[8]), .S(int_route_v[7]) ,.Q(int_resp_v[1]));
	MUX21X1 U24(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[9]), .S(int_route_v[7]) ,.Q(int_resp_v[2]));

	MUX21X1 U444(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[11]) ,.Q(int_map_req_v[444]));
	MUX21X1 U445(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[11]) ,.Q(int_map_req_v[445]));
	MUX21X1 U446(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[11]) ,.Q(int_map_req_v[446]));
	MUX21X1 U447(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[11]) ,.Q(int_map_req_v[447]));
	MUX21X1 U448(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[11]) ,.Q(int_map_req_v[448]));
	MUX21X1 U449(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[11]) ,.Q(int_map_req_v[449]));
	MUX21X1 U450(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[11]) ,.Q(int_map_req_v[450]));
	MUX21X1 U451(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[11]) ,.Q(int_map_req_v[451]));
	MUX21X1 U452(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[11]) ,.Q(int_map_req_v[452]));
	MUX21X1 U453(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[11]) ,.Q(int_map_req_v[453]));
	MUX21X1 U454(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[11]) ,.Q(int_map_req_v[454]));
	MUX21X1 U455(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[11]) ,.Q(int_map_req_v[455]));
	MUX21X1 U456(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[11]) ,.Q(int_map_req_v[456]));
	MUX21X1 U457(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[11]) ,.Q(int_map_req_v[457]));
	MUX21X1 U458(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[11]) ,.Q(int_map_req_v[458]));
	MUX21X1 U459(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[11]) ,.Q(int_map_req_v[459]));
	MUX21X1 U460(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[11]) ,.Q(int_map_req_v[460]));
	MUX21X1 U461(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[11]) ,.Q(int_map_req_v[461]));
	MUX21X1 U462(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[11]) ,.Q(int_map_req_v[462]));
	MUX21X1 U463(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[11]) ,.Q(int_map_req_v[463]));
	MUX21X1 U464(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[11]) ,.Q(int_map_req_v[464]));
	MUX21X1 U465(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[11]) ,.Q(int_map_req_v[465]));
	MUX21X1 U466(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[11]) ,.Q(int_map_req_v[466]));
	MUX21X1 U467(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[11]) ,.Q(int_map_req_v[467]));
	MUX21X1 U468(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[11]) ,.Q(int_map_req_v[468]));
	MUX21X1 U469(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[11]) ,.Q(int_map_req_v[469]));
	MUX21X1 U470(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[11]) ,.Q(int_map_req_v[470]));
	MUX21X1 U471(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[11]) ,.Q(int_map_req_v[471]));
	MUX21X1 U472(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[11]) ,.Q(int_map_req_v[472]));
	MUX21X1 U473(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[11]) ,.Q(int_map_req_v[473]));
	MUX21X1 U474(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[11]) ,.Q(int_map_req_v[474]));
	MUX21X1 U475(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[11]) ,.Q(int_map_req_v[475]));
	MUX21X1 U476(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[11]) ,.Q(int_map_req_v[476]));
	MUX21X1 U477(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[11]) ,.Q(int_map_req_v[477]));
	MUX21X1 U478(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[11]) ,.Q(int_map_req_v[478]));
	MUX21X1 U479(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[11]) ,.Q(int_map_req_v[479]));
	MUX21X1 U480(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[11]) ,.Q(int_map_req_v[480]));
	MUX21X1 U481(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[6]) ,.Q(int_map_req_v[481]));
	MUX21X1 U482(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[6]) ,.Q(int_map_req_v[482]));
	MUX21X1 U483(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[6]) ,.Q(int_map_req_v[483]));
	MUX21X1 U484(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[6]) ,.Q(int_map_req_v[484]));
	MUX21X1 U485(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[6]) ,.Q(int_map_req_v[485]));
	MUX21X1 U486(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[6]) ,.Q(int_map_req_v[486]));
	MUX21X1 U487(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[6]) ,.Q(int_map_req_v[487]));
	MUX21X1 U488(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[6]) ,.Q(int_map_req_v[488]));
	MUX21X1 U489(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[6]) ,.Q(int_map_req_v[489]));
	MUX21X1 U490(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[6]) ,.Q(int_map_req_v[490]));
	MUX21X1 U491(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[6]) ,.Q(int_map_req_v[491]));
	MUX21X1 U492(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[6]) ,.Q(int_map_req_v[492]));
	MUX21X1 U493(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[6]) ,.Q(int_map_req_v[493]));
	MUX21X1 U494(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[6]) ,.Q(int_map_req_v[494]));
	MUX21X1 U495(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[6]) ,.Q(int_map_req_v[495]));
	MUX21X1 U496(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[6]) ,.Q(int_map_req_v[496]));
	MUX21X1 U497(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[6]) ,.Q(int_map_req_v[497]));
	MUX21X1 U498(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[6]) ,.Q(int_map_req_v[498]));
	MUX21X1 U499(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[6]) ,.Q(int_map_req_v[499]));
	MUX21X1 U500(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[6]) ,.Q(int_map_req_v[500]));
	MUX21X1 U501(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[6]) ,.Q(int_map_req_v[501]));
	MUX21X1 U502(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[6]) ,.Q(int_map_req_v[502]));
	MUX21X1 U503(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[6]) ,.Q(int_map_req_v[503]));
	MUX21X1 U504(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[6]) ,.Q(int_map_req_v[504]));
	MUX21X1 U505(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[6]) ,.Q(int_map_req_v[505]));
	MUX21X1 U506(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[6]) ,.Q(int_map_req_v[506]));
	MUX21X1 U507(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[6]) ,.Q(int_map_req_v[507]));
	MUX21X1 U508(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[6]) ,.Q(int_map_req_v[508]));
	MUX21X1 U509(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[6]) ,.Q(int_map_req_v[509]));
	MUX21X1 U510(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[6]) ,.Q(int_map_req_v[510]));
	MUX21X1 U511(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[6]) ,.Q(int_map_req_v[511]));
	MUX21X1 U512(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[6]) ,.Q(int_map_req_v[512]));
	MUX21X1 U513(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[6]) ,.Q(int_map_req_v[513]));
	MUX21X1 U514(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[6]) ,.Q(int_map_req_v[514]));
	MUX21X1 U515(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[6]) ,.Q(int_map_req_v[515]));
	MUX21X1 U516(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[6]) ,.Q(int_map_req_v[516]));
	MUX21X1 U517(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[6]) ,.Q(int_map_req_v[517]));
	MUX21X1 U518(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[1]) ,.Q(int_map_req_v[518]));
	MUX21X1 U519(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[1]) ,.Q(int_map_req_v[519]));
	MUX21X1 U520(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[1]) ,.Q(int_map_req_v[520]));
	MUX21X1 U521(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[1]) ,.Q(int_map_req_v[521]));
	MUX21X1 U522(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[1]) ,.Q(int_map_req_v[522]));
	MUX21X1 U523(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[1]) ,.Q(int_map_req_v[523]));
	MUX21X1 U524(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[1]) ,.Q(int_map_req_v[524]));
	MUX21X1 U525(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[1]) ,.Q(int_map_req_v[525]));
	MUX21X1 U526(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[1]) ,.Q(int_map_req_v[526]));
	MUX21X1 U527(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[1]) ,.Q(int_map_req_v[527]));
	MUX21X1 U528(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[1]) ,.Q(int_map_req_v[528]));
	MUX21X1 U529(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[1]) ,.Q(int_map_req_v[529]));
	MUX21X1 U530(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[1]) ,.Q(int_map_req_v[530]));
	MUX21X1 U531(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[1]) ,.Q(int_map_req_v[531]));
	MUX21X1 U532(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[1]) ,.Q(int_map_req_v[532]));
	MUX21X1 U533(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[1]) ,.Q(int_map_req_v[533]));
	MUX21X1 U534(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[1]) ,.Q(int_map_req_v[534]));
	MUX21X1 U535(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[1]) ,.Q(int_map_req_v[535]));
	MUX21X1 U536(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[1]) ,.Q(int_map_req_v[536]));
	MUX21X1 U537(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[1]) ,.Q(int_map_req_v[537]));
	MUX21X1 U538(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[1]) ,.Q(int_map_req_v[538]));
	MUX21X1 U539(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[1]) ,.Q(int_map_req_v[539]));
	MUX21X1 U540(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[1]) ,.Q(int_map_req_v[540]));
	MUX21X1 U541(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[1]) ,.Q(int_map_req_v[541]));
	MUX21X1 U542(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[1]) ,.Q(int_map_req_v[542]));
	MUX21X1 U543(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[1]) ,.Q(int_map_req_v[543]));
	MUX21X1 U544(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[1]) ,.Q(int_map_req_v[544]));
	MUX21X1 U545(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[1]) ,.Q(int_map_req_v[545]));
	MUX21X1 U546(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[1]) ,.Q(int_map_req_v[546]));
	MUX21X1 U547(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[1]) ,.Q(int_map_req_v[547]));
	MUX21X1 U548(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[1]) ,.Q(int_map_req_v[548]));
	MUX21X1 U549(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[1]) ,.Q(int_map_req_v[549]));
	MUX21X1 U550(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[1]) ,.Q(int_map_req_v[550]));
	MUX21X1 U551(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[1]) ,.Q(int_map_req_v[551]));
	MUX21X1 U552(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[1]) ,.Q(int_map_req_v[552]));
	MUX21X1 U553(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[1]) ,.Q(int_map_req_v[553]));
	MUX21X1 U554(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[1]) ,.Q(int_map_req_v[554]));
	MUX21X1 U555(.IN1(1'sb0), .IN2(int_req_v[148]), .S(int_route_v[21]) ,.Q(int_map_req_v[555]));
	MUX21X1 U556(.IN1(1'sb0), .IN2(int_req_v[149]), .S(int_route_v[21]) ,.Q(int_map_req_v[556]));
	MUX21X1 U557(.IN1(1'sb0), .IN2(int_req_v[150]), .S(int_route_v[21]) ,.Q(int_map_req_v[557]));
	MUX21X1 U558(.IN1(1'sb0), .IN2(int_req_v[151]), .S(int_route_v[21]) ,.Q(int_map_req_v[558]));
	MUX21X1 U559(.IN1(1'sb0), .IN2(int_req_v[152]), .S(int_route_v[21]) ,.Q(int_map_req_v[559]));
	MUX21X1 U560(.IN1(1'sb0), .IN2(int_req_v[153]), .S(int_route_v[21]) ,.Q(int_map_req_v[560]));
	MUX21X1 U561(.IN1(1'sb0), .IN2(int_req_v[154]), .S(int_route_v[21]) ,.Q(int_map_req_v[561]));
	MUX21X1 U562(.IN1(1'sb0), .IN2(int_req_v[155]), .S(int_route_v[21]) ,.Q(int_map_req_v[562]));
	MUX21X1 U563(.IN1(1'sb0), .IN2(int_req_v[156]), .S(int_route_v[21]) ,.Q(int_map_req_v[563]));
	MUX21X1 U564(.IN1(1'sb0), .IN2(int_req_v[157]), .S(int_route_v[21]) ,.Q(int_map_req_v[564]));
	MUX21X1 U565(.IN1(1'sb0), .IN2(int_req_v[158]), .S(int_route_v[21]) ,.Q(int_map_req_v[565]));
	MUX21X1 U566(.IN1(1'sb0), .IN2(int_req_v[159]), .S(int_route_v[21]) ,.Q(int_map_req_v[566]));
	MUX21X1 U567(.IN1(1'sb0), .IN2(int_req_v[160]), .S(int_route_v[21]) ,.Q(int_map_req_v[567]));
	MUX21X1 U568(.IN1(1'sb0), .IN2(int_req_v[161]), .S(int_route_v[21]) ,.Q(int_map_req_v[568]));
	MUX21X1 U569(.IN1(1'sb0), .IN2(int_req_v[162]), .S(int_route_v[21]) ,.Q(int_map_req_v[569]));
	MUX21X1 U570(.IN1(1'sb0), .IN2(int_req_v[163]), .S(int_route_v[21]) ,.Q(int_map_req_v[570]));
	MUX21X1 U571(.IN1(1'sb0), .IN2(int_req_v[164]), .S(int_route_v[21]) ,.Q(int_map_req_v[571]));
	MUX21X1 U572(.IN1(1'sb0), .IN2(int_req_v[165]), .S(int_route_v[21]) ,.Q(int_map_req_v[572]));
	MUX21X1 U573(.IN1(1'sb0), .IN2(int_req_v[166]), .S(int_route_v[21]) ,.Q(int_map_req_v[573]));
	MUX21X1 U574(.IN1(1'sb0), .IN2(int_req_v[167]), .S(int_route_v[21]) ,.Q(int_map_req_v[574]));
	MUX21X1 U575(.IN1(1'sb0), .IN2(int_req_v[168]), .S(int_route_v[21]) ,.Q(int_map_req_v[575]));
	MUX21X1 U576(.IN1(1'sb0), .IN2(int_req_v[169]), .S(int_route_v[21]) ,.Q(int_map_req_v[576]));
	MUX21X1 U577(.IN1(1'sb0), .IN2(int_req_v[170]), .S(int_route_v[21]) ,.Q(int_map_req_v[577]));
	MUX21X1 U578(.IN1(1'sb0), .IN2(int_req_v[171]), .S(int_route_v[21]) ,.Q(int_map_req_v[578]));
	MUX21X1 U579(.IN1(1'sb0), .IN2(int_req_v[172]), .S(int_route_v[21]) ,.Q(int_map_req_v[579]));
	MUX21X1 U580(.IN1(1'sb0), .IN2(int_req_v[173]), .S(int_route_v[21]) ,.Q(int_map_req_v[580]));
	MUX21X1 U581(.IN1(1'sb0), .IN2(int_req_v[174]), .S(int_route_v[21]) ,.Q(int_map_req_v[581]));
	MUX21X1 U582(.IN1(1'sb0), .IN2(int_req_v[175]), .S(int_route_v[21]) ,.Q(int_map_req_v[582]));
	MUX21X1 U583(.IN1(1'sb0), .IN2(int_req_v[176]), .S(int_route_v[21]) ,.Q(int_map_req_v[583]));
	MUX21X1 U584(.IN1(1'sb0), .IN2(int_req_v[177]), .S(int_route_v[21]) ,.Q(int_map_req_v[584]));
	MUX21X1 U585(.IN1(1'sb0), .IN2(int_req_v[178]), .S(int_route_v[21]) ,.Q(int_map_req_v[585]));
	MUX21X1 U586(.IN1(1'sb0), .IN2(int_req_v[179]), .S(int_route_v[21]) ,.Q(int_map_req_v[586]));
	MUX21X1 U587(.IN1(1'sb0), .IN2(int_req_v[180]), .S(int_route_v[21]) ,.Q(int_map_req_v[587]));
	MUX21X1 U588(.IN1(1'sb0), .IN2(int_req_v[181]), .S(int_route_v[21]) ,.Q(int_map_req_v[588]));
	MUX21X1 U589(.IN1(1'sb0), .IN2(int_req_v[182]), .S(int_route_v[21]) ,.Q(int_map_req_v[589]));
	MUX21X1 U590(.IN1(1'sb0), .IN2(int_req_v[183]), .S(int_route_v[21]) ,.Q(int_map_req_v[590]));
	MUX21X1 U591(.IN1(1'sb0), .IN2(int_req_v[184]), .S(int_route_v[21]) ,.Q(int_map_req_v[591]));
	MUX21X1 U25(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[15]), .S(int_route_v[21]) ,.Q(int_resp_v[4]));
	MUX21X1 U26(.IN1(int_resp_v[5]), .IN2(int_map_resp_v[16]), .S(int_route_v[21]) ,.Q(int_resp_v[5]));
	MUX21X1 U27(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[14]), .S(int_route_v[1]) ,.Q(int_resp_v[0]));
	MUX21X1 U28(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[15]), .S(int_route_v[1]) ,.Q(int_resp_v[1]));
	MUX21X1 U29(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[13]), .S(int_route_v[6]) ,.Q(int_resp_v[1]));
	MUX21X1 U30(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[14]), .S(int_route_v[6]) ,.Q(int_resp_v[2]));
	MUX21X1 U31(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[12]), .S(int_route_v[11]) ,.Q(int_resp_v[2]));
	MUX21X1 U32(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[13]), .S(int_route_v[11]) ,.Q(int_resp_v[3]));



	MUX21X1 U592(.IN1(1'sb0), .IN2(int_req_v[111]), .S(int_route_v[15]) ,.Q(int_map_req_v[592]));
	MUX21X1 U593(.IN1(1'sb0), .IN2(int_req_v[112]), .S(int_route_v[15]) ,.Q(int_map_req_v[593]));
	MUX21X1 U594(.IN1(1'sb0), .IN2(int_req_v[113]), .S(int_route_v[15]) ,.Q(int_map_req_v[594]));
	MUX21X1 U595(.IN1(1'sb0), .IN2(int_req_v[114]), .S(int_route_v[15]) ,.Q(int_map_req_v[595]));
	MUX21X1 U596(.IN1(1'sb0), .IN2(int_req_v[115]), .S(int_route_v[15]) ,.Q(int_map_req_v[596]));
	MUX21X1 U597(.IN1(1'sb0), .IN2(int_req_v[116]), .S(int_route_v[15]) ,.Q(int_map_req_v[597]));
	MUX21X1 U598(.IN1(1'sb0), .IN2(int_req_v[117]), .S(int_route_v[15]) ,.Q(int_map_req_v[598]));
	MUX21X1 U599(.IN1(1'sb0), .IN2(int_req_v[118]), .S(int_route_v[15]) ,.Q(int_map_req_v[599]));
	MUX21X1 U600(.IN1(1'sb0), .IN2(int_req_v[119]), .S(int_route_v[15]) ,.Q(int_map_req_v[600]));
	MUX21X1 U601(.IN1(1'sb0), .IN2(int_req_v[120]), .S(int_route_v[15]) ,.Q(int_map_req_v[601]));
	MUX21X1 U602(.IN1(1'sb0), .IN2(int_req_v[121]), .S(int_route_v[15]) ,.Q(int_map_req_v[602]));
	MUX21X1 U603(.IN1(1'sb0), .IN2(int_req_v[122]), .S(int_route_v[15]) ,.Q(int_map_req_v[603]));
	MUX21X1 U604(.IN1(1'sb0), .IN2(int_req_v[123]), .S(int_route_v[15]) ,.Q(int_map_req_v[604]));
	MUX21X1 U605(.IN1(1'sb0), .IN2(int_req_v[124]), .S(int_route_v[15]) ,.Q(int_map_req_v[605]));
	MUX21X1 U606(.IN1(1'sb0), .IN2(int_req_v[125]), .S(int_route_v[15]) ,.Q(int_map_req_v[606]));
	MUX21X1 U607(.IN1(1'sb0), .IN2(int_req_v[126]), .S(int_route_v[15]) ,.Q(int_map_req_v[607]));
	MUX21X1 U608(.IN1(1'sb0), .IN2(int_req_v[127]), .S(int_route_v[15]) ,.Q(int_map_req_v[608]));
	MUX21X1 U609(.IN1(1'sb0), .IN2(int_req_v[128]), .S(int_route_v[15]) ,.Q(int_map_req_v[609]));
	MUX21X1 U610(.IN1(1'sb0), .IN2(int_req_v[129]), .S(int_route_v[15]) ,.Q(int_map_req_v[610]));
	MUX21X1 U611(.IN1(1'sb0), .IN2(int_req_v[130]), .S(int_route_v[15]) ,.Q(int_map_req_v[611]));
	MUX21X1 U612(.IN1(1'sb0), .IN2(int_req_v[131]), .S(int_route_v[15]) ,.Q(int_map_req_v[612]));
	MUX21X1 U613(.IN1(1'sb0), .IN2(int_req_v[132]), .S(int_route_v[15]) ,.Q(int_map_req_v[613]));
	MUX21X1 U614(.IN1(1'sb0), .IN2(int_req_v[133]), .S(int_route_v[15]) ,.Q(int_map_req_v[614]));
	MUX21X1 U615(.IN1(1'sb0), .IN2(int_req_v[134]), .S(int_route_v[15]) ,.Q(int_map_req_v[615]));
	MUX21X1 U616(.IN1(1'sb0), .IN2(int_req_v[135]), .S(int_route_v[15]) ,.Q(int_map_req_v[616]));
	MUX21X1 U617(.IN1(1'sb0), .IN2(int_req_v[136]), .S(int_route_v[15]) ,.Q(int_map_req_v[617]));
	MUX21X1 U618(.IN1(1'sb0), .IN2(int_req_v[137]), .S(int_route_v[15]) ,.Q(int_map_req_v[618]));
	MUX21X1 U619(.IN1(1'sb0), .IN2(int_req_v[138]), .S(int_route_v[15]) ,.Q(int_map_req_v[619]));
	MUX21X1 U620(.IN1(1'sb0), .IN2(int_req_v[139]), .S(int_route_v[15]) ,.Q(int_map_req_v[620]));
	MUX21X1 U621(.IN1(1'sb0), .IN2(int_req_v[140]), .S(int_route_v[15]) ,.Q(int_map_req_v[621]));
	MUX21X1 U622(.IN1(1'sb0), .IN2(int_req_v[141]), .S(int_route_v[15]) ,.Q(int_map_req_v[622]));
	MUX21X1 U623(.IN1(1'sb0), .IN2(int_req_v[142]), .S(int_route_v[15]) ,.Q(int_map_req_v[623]));
	MUX21X1 U624(.IN1(1'sb0), .IN2(int_req_v[143]), .S(int_route_v[15]) ,.Q(int_map_req_v[624]));
	MUX21X1 U625(.IN1(1'sb0), .IN2(int_req_v[144]), .S(int_route_v[15]) ,.Q(int_map_req_v[625]));
	MUX21X1 U626(.IN1(1'sb0), .IN2(int_req_v[145]), .S(int_route_v[15]) ,.Q(int_map_req_v[626]));
	MUX21X1 U627(.IN1(1'sb0), .IN2(int_req_v[146]), .S(int_route_v[15]) ,.Q(int_map_req_v[627]));
	MUX21X1 U628(.IN1(1'sb0), .IN2(int_req_v[147]), .S(int_route_v[15]) ,.Q(int_map_req_v[628]));
	MUX21X1 U629(.IN1(1'sb0), .IN2(int_req_v[74]), .S(int_route_v[10]) ,.Q(int_map_req_v[629]));
	MUX21X1 U630(.IN1(1'sb0), .IN2(int_req_v[75]), .S(int_route_v[10]) ,.Q(int_map_req_v[630]));
	MUX21X1 U631(.IN1(1'sb0), .IN2(int_req_v[76]), .S(int_route_v[10]) ,.Q(int_map_req_v[631]));
	MUX21X1 U632(.IN1(1'sb0), .IN2(int_req_v[77]), .S(int_route_v[10]) ,.Q(int_map_req_v[632]));
	MUX21X1 U633(.IN1(1'sb0), .IN2(int_req_v[78]), .S(int_route_v[10]) ,.Q(int_map_req_v[633]));
	MUX21X1 U634(.IN1(1'sb0), .IN2(int_req_v[79]), .S(int_route_v[10]) ,.Q(int_map_req_v[634]));
	MUX21X1 U635(.IN1(1'sb0), .IN2(int_req_v[80]), .S(int_route_v[10]) ,.Q(int_map_req_v[635]));
	MUX21X1 U636(.IN1(1'sb0), .IN2(int_req_v[81]), .S(int_route_v[10]) ,.Q(int_map_req_v[636]));
	MUX21X1 U637(.IN1(1'sb0), .IN2(int_req_v[82]), .S(int_route_v[10]) ,.Q(int_map_req_v[637]));
	MUX21X1 U638(.IN1(1'sb0), .IN2(int_req_v[83]), .S(int_route_v[10]) ,.Q(int_map_req_v[638]));
	MUX21X1 U639(.IN1(1'sb0), .IN2(int_req_v[84]), .S(int_route_v[10]) ,.Q(int_map_req_v[639]));
	MUX21X1 U640(.IN1(1'sb0), .IN2(int_req_v[85]), .S(int_route_v[10]) ,.Q(int_map_req_v[640]));
	MUX21X1 U641(.IN1(1'sb0), .IN2(int_req_v[86]), .S(int_route_v[10]) ,.Q(int_map_req_v[641]));
	MUX21X1 U642(.IN1(1'sb0), .IN2(int_req_v[87]), .S(int_route_v[10]) ,.Q(int_map_req_v[642]));
	MUX21X1 U643(.IN1(1'sb0), .IN2(int_req_v[88]), .S(int_route_v[10]) ,.Q(int_map_req_v[643]));
	MUX21X1 U644(.IN1(1'sb0), .IN2(int_req_v[89]), .S(int_route_v[10]) ,.Q(int_map_req_v[644]));
	MUX21X1 U645(.IN1(1'sb0), .IN2(int_req_v[90]), .S(int_route_v[10]) ,.Q(int_map_req_v[645]));
	MUX21X1 U646(.IN1(1'sb0), .IN2(int_req_v[91]), .S(int_route_v[10]) ,.Q(int_map_req_v[646]));
	MUX21X1 U647(.IN1(1'sb0), .IN2(int_req_v[92]), .S(int_route_v[10]) ,.Q(int_map_req_v[647]));
	MUX21X1 U648(.IN1(1'sb0), .IN2(int_req_v[93]), .S(int_route_v[10]) ,.Q(int_map_req_v[648]));
	MUX21X1 U649(.IN1(1'sb0), .IN2(int_req_v[94]), .S(int_route_v[10]) ,.Q(int_map_req_v[649]));
	MUX21X1 U650(.IN1(1'sb0), .IN2(int_req_v[95]), .S(int_route_v[10]) ,.Q(int_map_req_v[650]));
	MUX21X1 U651(.IN1(1'sb0), .IN2(int_req_v[96]), .S(int_route_v[10]) ,.Q(int_map_req_v[651]));
	MUX21X1 U652(.IN1(1'sb0), .IN2(int_req_v[97]), .S(int_route_v[10]) ,.Q(int_map_req_v[652]));
	MUX21X1 U653(.IN1(1'sb0), .IN2(int_req_v[98]), .S(int_route_v[10]) ,.Q(int_map_req_v[653]));
	MUX21X1 U654(.IN1(1'sb0), .IN2(int_req_v[99]), .S(int_route_v[10]) ,.Q(int_map_req_v[654]));
	MUX21X1 U655(.IN1(1'sb0), .IN2(int_req_v[100]), .S(int_route_v[10]) ,.Q(int_map_req_v[655]));
	MUX21X1 U656(.IN1(1'sb0), .IN2(int_req_v[101]), .S(int_route_v[10]) ,.Q(int_map_req_v[656]));
	MUX21X1 U657(.IN1(1'sb0), .IN2(int_req_v[102]), .S(int_route_v[10]) ,.Q(int_map_req_v[657]));
	MUX21X1 U658(.IN1(1'sb0), .IN2(int_req_v[103]), .S(int_route_v[10]) ,.Q(int_map_req_v[658]));
	MUX21X1 U659(.IN1(1'sb0), .IN2(int_req_v[104]), .S(int_route_v[10]) ,.Q(int_map_req_v[659]));
	MUX21X1 U660(.IN1(1'sb0), .IN2(int_req_v[105]), .S(int_route_v[10]) ,.Q(int_map_req_v[660]));
	MUX21X1 U661(.IN1(1'sb0), .IN2(int_req_v[106]), .S(int_route_v[10]) ,.Q(int_map_req_v[661]));
	MUX21X1 U662(.IN1(1'sb0), .IN2(int_req_v[107]), .S(int_route_v[10]) ,.Q(int_map_req_v[662]));
	MUX21X1 U663(.IN1(1'sb0), .IN2(int_req_v[108]), .S(int_route_v[10]) ,.Q(int_map_req_v[663]));
	MUX21X1 U664(.IN1(1'sb0), .IN2(int_req_v[109]), .S(int_route_v[10]) ,.Q(int_map_req_v[664]));
	MUX21X1 U665(.IN1(1'sb0), .IN2(int_req_v[110]), .S(int_route_v[10]) ,.Q(int_map_req_v[665]));
	MUX21X1 U666(.IN1(1'sb0), .IN2(int_req_v[37]), .S(int_route_v[5]) ,.Q(int_map_req_v[666]));
	MUX21X1 U667(.IN1(1'sb0), .IN2(int_req_v[38]), .S(int_route_v[5]) ,.Q(int_map_req_v[667]));
	MUX21X1 U668(.IN1(1'sb0), .IN2(int_req_v[39]), .S(int_route_v[5]) ,.Q(int_map_req_v[668]));
	MUX21X1 U669(.IN1(1'sb0), .IN2(int_req_v[40]), .S(int_route_v[5]) ,.Q(int_map_req_v[669]));
	MUX21X1 U670(.IN1(1'sb0), .IN2(int_req_v[41]), .S(int_route_v[5]) ,.Q(int_map_req_v[670]));
	MUX21X1 U671(.IN1(1'sb0), .IN2(int_req_v[42]), .S(int_route_v[5]) ,.Q(int_map_req_v[671]));
	MUX21X1 U672(.IN1(1'sb0), .IN2(int_req_v[43]), .S(int_route_v[5]) ,.Q(int_map_req_v[672]));
	MUX21X1 U673(.IN1(1'sb0), .IN2(int_req_v[44]), .S(int_route_v[5]) ,.Q(int_map_req_v[673]));
	MUX21X1 U674(.IN1(1'sb0), .IN2(int_req_v[45]), .S(int_route_v[5]) ,.Q(int_map_req_v[674]));
	MUX21X1 U675(.IN1(1'sb0), .IN2(int_req_v[46]), .S(int_route_v[5]) ,.Q(int_map_req_v[675]));
	MUX21X1 U676(.IN1(1'sb0), .IN2(int_req_v[47]), .S(int_route_v[5]) ,.Q(int_map_req_v[676]));
	MUX21X1 U677(.IN1(1'sb0), .IN2(int_req_v[48]), .S(int_route_v[5]) ,.Q(int_map_req_v[677]));
	MUX21X1 U678(.IN1(1'sb0), .IN2(int_req_v[49]), .S(int_route_v[5]) ,.Q(int_map_req_v[678]));
	MUX21X1 U679(.IN1(1'sb0), .IN2(int_req_v[50]), .S(int_route_v[5]) ,.Q(int_map_req_v[679]));
	MUX21X1 U680(.IN1(1'sb0), .IN2(int_req_v[51]), .S(int_route_v[5]) ,.Q(int_map_req_v[680]));
	MUX21X1 U681(.IN1(1'sb0), .IN2(int_req_v[52]), .S(int_route_v[5]) ,.Q(int_map_req_v[681]));
	MUX21X1 U682(.IN1(1'sb0), .IN2(int_req_v[53]), .S(int_route_v[5]) ,.Q(int_map_req_v[682]));
	MUX21X1 U683(.IN1(1'sb0), .IN2(int_req_v[54]), .S(int_route_v[5]) ,.Q(int_map_req_v[683]));
	MUX21X1 U684(.IN1(1'sb0), .IN2(int_req_v[55]), .S(int_route_v[5]) ,.Q(int_map_req_v[684]));
	MUX21X1 U685(.IN1(1'sb0), .IN2(int_req_v[56]), .S(int_route_v[5]) ,.Q(int_map_req_v[685]));
	MUX21X1 U686(.IN1(1'sb0), .IN2(int_req_v[57]), .S(int_route_v[5]) ,.Q(int_map_req_v[686]));
	MUX21X1 U687(.IN1(1'sb0), .IN2(int_req_v[58]), .S(int_route_v[5]) ,.Q(int_map_req_v[687]));
	MUX21X1 U688(.IN1(1'sb0), .IN2(int_req_v[59]), .S(int_route_v[5]) ,.Q(int_map_req_v[688]));
	MUX21X1 U689(.IN1(1'sb0), .IN2(int_req_v[60]), .S(int_route_v[5]) ,.Q(int_map_req_v[689]));
	MUX21X1 U690(.IN1(1'sb0), .IN2(int_req_v[61]), .S(int_route_v[5]) ,.Q(int_map_req_v[690]));
	MUX21X1 U691(.IN1(1'sb0), .IN2(int_req_v[62]), .S(int_route_v[5]) ,.Q(int_map_req_v[691]));
	MUX21X1 U692(.IN1(1'sb0), .IN2(int_req_v[63]), .S(int_route_v[5]) ,.Q(int_map_req_v[692]));
	MUX21X1 U693(.IN1(1'sb0), .IN2(int_req_v[64]), .S(int_route_v[5]) ,.Q(int_map_req_v[693]));
	MUX21X1 U694(.IN1(1'sb0), .IN2(int_req_v[65]), .S(int_route_v[5]) ,.Q(int_map_req_v[694]));
	MUX21X1 U695(.IN1(1'sb0), .IN2(int_req_v[66]), .S(int_route_v[5]) ,.Q(int_map_req_v[695]));
	MUX21X1 U696(.IN1(1'sb0), .IN2(int_req_v[67]), .S(int_route_v[5]) ,.Q(int_map_req_v[696]));
	MUX21X1 U697(.IN1(1'sb0), .IN2(int_req_v[68]), .S(int_route_v[5]) ,.Q(int_map_req_v[697]));
	MUX21X1 U698(.IN1(1'sb0), .IN2(int_req_v[69]), .S(int_route_v[5]) ,.Q(int_map_req_v[698]));
	MUX21X1 U699(.IN1(1'sb0), .IN2(int_req_v[70]), .S(int_route_v[5]) ,.Q(int_map_req_v[699]));
	MUX21X1 U700(.IN1(1'sb0), .IN2(int_req_v[71]), .S(int_route_v[5]) ,.Q(int_map_req_v[700]));
	MUX21X1 U701(.IN1(1'sb0), .IN2(int_req_v[72]), .S(int_route_v[5]) ,.Q(int_map_req_v[701]));
	MUX21X1 U702(.IN1(1'sb0), .IN2(int_req_v[73]), .S(int_route_v[5]) ,.Q(int_map_req_v[702]));
	MUX21X1 U703(.IN1(1'sb0), .IN2(int_req_v[0]), .S(int_route_v[0]) ,.Q(int_map_req_v[703]));
	MUX21X1 U704(.IN1(1'sb0), .IN2(int_req_v[1]), .S(int_route_v[0]) ,.Q(int_map_req_v[704]));
	MUX21X1 U705(.IN1(1'sb0), .IN2(int_req_v[2]), .S(int_route_v[0]) ,.Q(int_map_req_v[705]));
	MUX21X1 U706(.IN1(1'sb0), .IN2(int_req_v[3]), .S(int_route_v[0]) ,.Q(int_map_req_v[706]));
	MUX21X1 U707(.IN1(1'sb0), .IN2(int_req_v[4]), .S(int_route_v[0]) ,.Q(int_map_req_v[707]));
	MUX21X1 U708(.IN1(1'sb0), .IN2(int_req_v[5]), .S(int_route_v[0]) ,.Q(int_map_req_v[708]));
	MUX21X1 U709(.IN1(1'sb0), .IN2(int_req_v[6]), .S(int_route_v[0]) ,.Q(int_map_req_v[709]));
	MUX21X1 U710(.IN1(1'sb0), .IN2(int_req_v[7]), .S(int_route_v[0]) ,.Q(int_map_req_v[710]));
	MUX21X1 U711(.IN1(1'sb0), .IN2(int_req_v[8]), .S(int_route_v[0]) ,.Q(int_map_req_v[711]));
	MUX21X1 U712(.IN1(1'sb0), .IN2(int_req_v[9]), .S(int_route_v[0]) ,.Q(int_map_req_v[712]));
	MUX21X1 U713(.IN1(1'sb0), .IN2(int_req_v[10]), .S(int_route_v[0]) ,.Q(int_map_req_v[713]));
	MUX21X1 U714(.IN1(1'sb0), .IN2(int_req_v[11]), .S(int_route_v[0]) ,.Q(int_map_req_v[714]));
	MUX21X1 U715(.IN1(1'sb0), .IN2(int_req_v[12]), .S(int_route_v[0]) ,.Q(int_map_req_v[715]));
	MUX21X1 U716(.IN1(1'sb0), .IN2(int_req_v[13]), .S(int_route_v[0]) ,.Q(int_map_req_v[716]));
	MUX21X1 U717(.IN1(1'sb0), .IN2(int_req_v[14]), .S(int_route_v[0]) ,.Q(int_map_req_v[717]));
	MUX21X1 U718(.IN1(1'sb0), .IN2(int_req_v[15]), .S(int_route_v[0]) ,.Q(int_map_req_v[718]));
	MUX21X1 U719(.IN1(1'sb0), .IN2(int_req_v[16]), .S(int_route_v[0]) ,.Q(int_map_req_v[719]));
	MUX21X1 U720(.IN1(1'sb0), .IN2(int_req_v[17]), .S(int_route_v[0]) ,.Q(int_map_req_v[720]));
	MUX21X1 U721(.IN1(1'sb0), .IN2(int_req_v[18]), .S(int_route_v[0]) ,.Q(int_map_req_v[721]));
	MUX21X1 U722(.IN1(1'sb0), .IN2(int_req_v[19]), .S(int_route_v[0]) ,.Q(int_map_req_v[722]));
	MUX21X1 U723(.IN1(1'sb0), .IN2(int_req_v[20]), .S(int_route_v[0]) ,.Q(int_map_req_v[723]));
	MUX21X1 U724(.IN1(1'sb0), .IN2(int_req_v[21]), .S(int_route_v[0]) ,.Q(int_map_req_v[724]));
	MUX21X1 U725(.IN1(1'sb0), .IN2(int_req_v[22]), .S(int_route_v[0]) ,.Q(int_map_req_v[725]));
	MUX21X1 U726(.IN1(1'sb0), .IN2(int_req_v[23]), .S(int_route_v[0]) ,.Q(int_map_req_v[726]));
	MUX21X1 U727(.IN1(1'sb0), .IN2(int_req_v[24]), .S(int_route_v[0]) ,.Q(int_map_req_v[727]));
	MUX21X1 U728(.IN1(1'sb0), .IN2(int_req_v[25]), .S(int_route_v[0]) ,.Q(int_map_req_v[728]));
	MUX21X1 U729(.IN1(1'sb0), .IN2(int_req_v[26]), .S(int_route_v[0]) ,.Q(int_map_req_v[729]));
	MUX21X1 U730(.IN1(1'sb0), .IN2(int_req_v[27]), .S(int_route_v[0]) ,.Q(int_map_req_v[730]));
	MUX21X1 U731(.IN1(1'sb0), .IN2(int_req_v[28]), .S(int_route_v[0]) ,.Q(int_map_req_v[731]));
	MUX21X1 U732(.IN1(1'sb0), .IN2(int_req_v[29]), .S(int_route_v[0]) ,.Q(int_map_req_v[732]));
	MUX21X1 U733(.IN1(1'sb0), .IN2(int_req_v[30]), .S(int_route_v[0]) ,.Q(int_map_req_v[733]));
	MUX21X1 U734(.IN1(1'sb0), .IN2(int_req_v[31]), .S(int_route_v[0]) ,.Q(int_map_req_v[734]));
	MUX21X1 U735(.IN1(1'sb0), .IN2(int_req_v[32]), .S(int_route_v[0]) ,.Q(int_map_req_v[735]));
	MUX21X1 U736(.IN1(1'sb0), .IN2(int_req_v[33]), .S(int_route_v[0]) ,.Q(int_map_req_v[736]));
	MUX21X1 U737(.IN1(1'sb0), .IN2(int_req_v[34]), .S(int_route_v[0]) ,.Q(int_map_req_v[737]));
	MUX21X1 U738(.IN1(1'sb0), .IN2(int_req_v[35]), .S(int_route_v[0]) ,.Q(int_map_req_v[738]));
	MUX21X1 U739(.IN1(1'sb0), .IN2(int_req_v[36]), .S(int_route_v[0]) ,.Q(int_map_req_v[739]));
	MUX21X1 U33(.IN1(int_resp_v[0]), .IN2(int_map_resp_v[19]), .S(int_route_v[0]) ,.Q(int_resp_v[0]));
	MUX21X1 U34(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[20]), .S(int_route_v[0]) ,.Q(int_resp_v[1]));
	MUX21X1 U35(.IN1(int_resp_v[1]), .IN2(int_map_resp_v[18]), .S(int_route_v[5]) ,.Q(int_resp_v[1]));
	MUX21X1 U36(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[19]), .S(int_route_v[5]) ,.Q(int_resp_v[2]));
	MUX21X1 U37(.IN1(int_resp_v[2]), .IN2(int_map_resp_v[17]), .S(int_route_v[10]) ,.Q(int_resp_v[2]));
	MUX21X1 U38(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[18]), .S(int_route_v[10]) ,.Q(int_resp_v[3]));
	MUX21X1 U39(.IN1(int_resp_v[3]), .IN2(int_map_resp_v[16]), .S(int_route_v[15]) ,.Q(int_resp_v[3]));
	MUX21X1 U40(.IN1(int_resp_v[4]), .IN2(int_map_resp_v[17]), .S(int_route_v[15]) ,.Q(int_resp_v[4]));
